
`timescale 1ns/1ps
module mem_bram #(
    parameter ADDR_WIDTH = 10,		//地址宽度
    parameter DATA_WIDTH = 128		//数据宽度
)(
    input                   clk,   // Clock
    input [ADDR_WIDTH-1:0]  raddr,  // Address
    input [ADDR_WIDTH-1:0]  waddr,  // Address
    input [DATA_WIDTH-1:0]  din,   // Data Input
    input                   we,    // Write Enable
    output [DATA_WIDTH-1:0] dout   // Data Output
); 
    reg [ADDR_WIDTH-1:0] addr_r;  // Address Register
    reg [DATA_WIDTH-1:0] ram [0:(1 << ADDR_WIDTH)-1];
    integer i;
    initial begin
        ram[0][31:0] = 32'd726190305;
        ram[0][63:32] = 32'd855531051;
        ram[0][95:64] = 32'd2127818576;
        ram[0][127:96] = 32'd2710397198;
        ram[1][31:0] = 32'd919744787;
        ram[1][63:32] = 32'd1473416459;
        ram[1][95:64] = 32'd469065942;
        ram[1][127:96] = 32'd2410401329;
        ram[2][31:0] = 32'd1070477180;
        ram[2][63:32] = 32'd536276757;
        ram[2][95:64] = 32'd4272705751;
        ram[2][127:96] = 32'd1048550729;
        ram[3][31:0] = 32'd1981417174;
        ram[3][63:32] = 32'd467742172;
        ram[3][95:64] = 32'd3538414074;
        ram[3][127:96] = 32'd87988345;
        ram[4][31:0] = 32'd3931434522;
        ram[4][63:32] = 32'd3004992471;
        ram[4][95:64] = 32'd3664118966;
        ram[4][127:96] = 32'd2697384543;
        ram[5][31:0] = 32'd3947163269;
        ram[5][63:32] = 32'd789026206;
        ram[5][95:64] = 32'd2308919392;
        ram[5][127:96] = 32'd2328303965;
        ram[6][31:0] = 32'd3510174251;
        ram[6][63:32] = 32'd135025247;
        ram[6][95:64] = 32'd884555627;
        ram[6][127:96] = 32'd56674262;
        ram[7][31:0] = 32'd3998150063;
        ram[7][63:32] = 32'd4050089466;
        ram[7][95:64] = 32'd561337608;
        ram[7][127:96] = 32'd2160288399;
        ram[8][31:0] = 32'd2185218372;
        ram[8][63:32] = 32'd3281604318;
        ram[8][95:64] = 32'd3632025959;
        ram[8][127:96] = 32'd3955127962;
        ram[9][31:0] = 32'd3896309806;
        ram[9][63:32] = 32'd3905953463;
        ram[9][95:64] = 32'd1762764931;
        ram[9][127:96] = 32'd1468237573;
        ram[10][31:0] = 32'd3594722951;
        ram[10][63:32] = 32'd786275004;
        ram[10][95:64] = 32'd4096363574;
        ram[10][127:96] = 32'd3562471067;
        ram[11][31:0] = 32'd3885394360;
        ram[11][63:32] = 32'd720913470;
        ram[11][95:64] = 32'd2323962822;
        ram[11][127:96] = 32'd658713850;
        ram[12][31:0] = 32'd3954156962;
        ram[12][63:32] = 32'd2053400777;
        ram[12][95:64] = 32'd2548991497;
        ram[12][127:96] = 32'd869359556;
        ram[13][31:0] = 32'd3694524907;
        ram[13][63:32] = 32'd1440417870;
        ram[13][95:64] = 32'd3762075597;
        ram[13][127:96] = 32'd812389879;
        ram[14][31:0] = 32'd897892176;
        ram[14][63:32] = 32'd2822047506;
        ram[14][95:64] = 32'd2365235314;
        ram[14][127:96] = 32'd1947913714;
        ram[15][31:0] = 32'd3343706505;
        ram[15][63:32] = 32'd3050866392;
        ram[15][95:64] = 32'd389109591;
        ram[15][127:96] = 32'd3604968536;
        ram[16][31:0] = 32'd1958157960;
        ram[16][63:32] = 32'd2483132969;
        ram[16][95:64] = 32'd1363225947;
        ram[16][127:96] = 32'd3709922740;
        ram[17][31:0] = 32'd780007243;
        ram[17][63:32] = 32'd445386276;
        ram[17][95:64] = 32'd2608166339;
        ram[17][127:96] = 32'd1938766220;
        ram[18][31:0] = 32'd1907660428;
        ram[18][63:32] = 32'd261290754;
        ram[18][95:64] = 32'd1838785218;
        ram[18][127:96] = 32'd2999248499;
        ram[19][31:0] = 32'd1148223066;
        ram[19][63:32] = 32'd57221148;
        ram[19][95:64] = 32'd3865815998;
        ram[19][127:96] = 32'd4243798425;
        ram[20][31:0] = 32'd3551938821;
        ram[20][63:32] = 32'd2361350250;
        ram[20][95:64] = 32'd2006336925;
        ram[20][127:96] = 32'd4027428377;
        ram[21][31:0] = 32'd2985065750;
        ram[21][63:32] = 32'd1348591937;
        ram[21][95:64] = 32'd2748145392;
        ram[21][127:96] = 32'd3337487982;
        ram[22][31:0] = 32'd1328154912;
        ram[22][63:32] = 32'd4216399496;
        ram[22][95:64] = 32'd684440951;
        ram[22][127:96] = 32'd4038100292;
        ram[23][31:0] = 32'd11431343;
        ram[23][63:32] = 32'd1418096384;
        ram[23][95:64] = 32'd4104930478;
        ram[23][127:96] = 32'd1692585587;
        ram[24][31:0] = 32'd767733627;
        ram[24][63:32] = 32'd62382029;
        ram[24][95:64] = 32'd611847547;
        ram[24][127:96] = 32'd962759878;
        ram[25][31:0] = 32'd3727187527;
        ram[25][63:32] = 32'd334015143;
        ram[25][95:64] = 32'd1684138397;
        ram[25][127:96] = 32'd3519285150;
        ram[26][31:0] = 32'd912554404;
        ram[26][63:32] = 32'd1192418195;
        ram[26][95:64] = 32'd1862545842;
        ram[26][127:96] = 32'd347323893;
        ram[27][31:0] = 32'd849662807;
        ram[27][63:32] = 32'd2687315092;
        ram[27][95:64] = 32'd1367281977;
        ram[27][127:96] = 32'd3145322533;
        ram[28][31:0] = 32'd1757482678;
        ram[28][63:32] = 32'd419860717;
        ram[28][95:64] = 32'd4093300057;
        ram[28][127:96] = 32'd2847575930;
        ram[29][31:0] = 32'd3290921176;
        ram[29][63:32] = 32'd2303502259;
        ram[29][95:64] = 32'd1346885424;
        ram[29][127:96] = 32'd3348202238;
        ram[30][31:0] = 32'd167610123;
        ram[30][63:32] = 32'd3447666879;
        ram[30][95:64] = 32'd2514466426;
        ram[30][127:96] = 32'd3166000446;
        ram[31][31:0] = 32'd72247830;
        ram[31][63:32] = 32'd682282384;
        ram[31][95:64] = 32'd3834634229;
        ram[31][127:96] = 32'd1143290961;
        ram[32][31:0] = 32'd2369463817;
        ram[32][63:32] = 32'd4027118416;
        ram[32][95:64] = 32'd939881898;
        ram[32][127:96] = 32'd3754095223;
        ram[33][31:0] = 32'd438108953;
        ram[33][63:32] = 32'd2160563348;
        ram[33][95:64] = 32'd3949239056;
        ram[33][127:96] = 32'd3089281077;
        ram[34][31:0] = 32'd933962107;
        ram[34][63:32] = 32'd4248940189;
        ram[34][95:64] = 32'd44804164;
        ram[34][127:96] = 32'd3271595497;
        ram[35][31:0] = 32'd484269002;
        ram[35][63:32] = 32'd2186149626;
        ram[35][95:64] = 32'd2263992737;
        ram[35][127:96] = 32'd4166209102;
        ram[36][31:0] = 32'd1720721755;
        ram[36][63:32] = 32'd1758650845;
        ram[36][95:64] = 32'd3243521201;
        ram[36][127:96] = 32'd3596274834;
        ram[37][31:0] = 32'd310279149;
        ram[37][63:32] = 32'd368857195;
        ram[37][95:64] = 32'd1520413704;
        ram[37][127:96] = 32'd4042063966;
        ram[38][31:0] = 32'd2706977723;
        ram[38][63:32] = 32'd2764886121;
        ram[38][95:64] = 32'd818530140;
        ram[38][127:96] = 32'd2168736915;
        ram[39][31:0] = 32'd3532809018;
        ram[39][63:32] = 32'd1886808711;
        ram[39][95:64] = 32'd3247124859;
        ram[39][127:96] = 32'd3848464431;
        ram[40][31:0] = 32'd205033297;
        ram[40][63:32] = 32'd2014229717;
        ram[40][95:64] = 32'd3110936348;
        ram[40][127:96] = 32'd4051124924;
        ram[41][31:0] = 32'd3104036377;
        ram[41][63:32] = 32'd190214731;
        ram[41][95:64] = 32'd3551362444;
        ram[41][127:96] = 32'd769142066;
        ram[42][31:0] = 32'd546345531;
        ram[42][63:32] = 32'd137499134;
        ram[42][95:64] = 32'd1650688480;
        ram[42][127:96] = 32'd2112141990;
        ram[43][31:0] = 32'd1681519392;
        ram[43][63:32] = 32'd2097875581;
        ram[43][95:64] = 32'd2644158774;
        ram[43][127:96] = 32'd2234447425;
        ram[44][31:0] = 32'd615319646;
        ram[44][63:32] = 32'd2905827243;
        ram[44][95:64] = 32'd3643073190;
        ram[44][127:96] = 32'd3882480974;
        ram[45][31:0] = 32'd1768002488;
        ram[45][63:32] = 32'd3711414204;
        ram[45][95:64] = 32'd3939676421;
        ram[45][127:96] = 32'd4082433942;
        ram[46][31:0] = 32'd3271992916;
        ram[46][63:32] = 32'd4056616662;
        ram[46][95:64] = 32'd3350085156;
        ram[46][127:96] = 32'd1241473016;
        ram[47][31:0] = 32'd3694204641;
        ram[47][63:32] = 32'd2413112707;
        ram[47][95:64] = 32'd3753406994;
        ram[47][127:96] = 32'd3616306016;
        ram[48][31:0] = 32'd1803940817;
        ram[48][63:32] = 32'd1827492103;
        ram[48][95:64] = 32'd2743985160;
        ram[48][127:96] = 32'd2074235098;
        ram[49][31:0] = 32'd1007003283;
        ram[49][63:32] = 32'd1022834255;
        ram[49][95:64] = 32'd3924284121;
        ram[49][127:96] = 32'd1949557997;
        ram[50][31:0] = 32'd187765645;
        ram[50][63:32] = 32'd2352154551;
        ram[50][95:64] = 32'd3541495957;
        ram[50][127:96] = 32'd1701074922;
        ram[51][31:0] = 32'd658105954;
        ram[51][63:32] = 32'd3083248378;
        ram[51][95:64] = 32'd2742135044;
        ram[51][127:96] = 32'd1009790862;
        ram[52][31:0] = 32'd881023582;
        ram[52][63:32] = 32'd3871168379;
        ram[52][95:64] = 32'd1795570751;
        ram[52][127:96] = 32'd3319553303;
        ram[53][31:0] = 32'd51944071;
        ram[53][63:32] = 32'd121162192;
        ram[53][95:64] = 32'd631424203;
        ram[53][127:96] = 32'd815101909;
        ram[54][31:0] = 32'd3992465811;
        ram[54][63:32] = 32'd2521597648;
        ram[54][95:64] = 32'd4290554056;
        ram[54][127:96] = 32'd1413986338;
        ram[55][31:0] = 32'd1246824563;
        ram[55][63:32] = 32'd2967623187;
        ram[55][95:64] = 32'd4085577484;
        ram[55][127:96] = 32'd3855190456;
        ram[56][31:0] = 32'd643551870;
        ram[56][63:32] = 32'd524980437;
        ram[56][95:64] = 32'd1741714033;
        ram[56][127:96] = 32'd480468405;
        ram[57][31:0] = 32'd1885599207;
        ram[57][63:32] = 32'd1480893710;
        ram[57][95:64] = 32'd2986628736;
        ram[57][127:96] = 32'd660798456;
        ram[58][31:0] = 32'd2070368912;
        ram[58][63:32] = 32'd2430721901;
        ram[58][95:64] = 32'd3326904585;
        ram[58][127:96] = 32'd3516786644;
        ram[59][31:0] = 32'd3976153366;
        ram[59][63:32] = 32'd1687762213;
        ram[59][95:64] = 32'd83366238;
        ram[59][127:96] = 32'd948945575;
        ram[60][31:0] = 32'd2608724663;
        ram[60][63:32] = 32'd1993840260;
        ram[60][95:64] = 32'd2171707476;
        ram[60][127:96] = 32'd1003754273;
        ram[61][31:0] = 32'd2164984734;
        ram[61][63:32] = 32'd1076761213;
        ram[61][95:64] = 32'd1264185063;
        ram[61][127:96] = 32'd4145441796;
        ram[62][31:0] = 32'd2470758762;
        ram[62][63:32] = 32'd4257985210;
        ram[62][95:64] = 32'd2354385756;
        ram[62][127:96] = 32'd3619119446;
        ram[63][31:0] = 32'd4126756018;
        ram[63][63:32] = 32'd3724959485;
        ram[63][95:64] = 32'd714648240;
        ram[63][127:96] = 32'd753719973;
        ram[64][31:0] = 32'd3872731299;
        ram[64][63:32] = 32'd2532794738;
        ram[64][95:64] = 32'd1832274105;
        ram[64][127:96] = 32'd1475111032;
        ram[65][31:0] = 32'd2709922654;
        ram[65][63:32] = 32'd3806634879;
        ram[65][95:64] = 32'd1218402663;
        ram[65][127:96] = 32'd1115477981;
        ram[66][31:0] = 32'd835312204;
        ram[66][63:32] = 32'd1680147033;
        ram[66][95:64] = 32'd2089647551;
        ram[66][127:96] = 32'd326083300;
        ram[67][31:0] = 32'd2027770644;
        ram[67][63:32] = 32'd478738172;
        ram[67][95:64] = 32'd3662961798;
        ram[67][127:96] = 32'd3753349860;
        ram[68][31:0] = 32'd3167753977;
        ram[68][63:32] = 32'd2277303350;
        ram[68][95:64] = 32'd3059293611;
        ram[68][127:96] = 32'd2980684711;
        ram[69][31:0] = 32'd3748482894;
        ram[69][63:32] = 32'd2128154341;
        ram[69][95:64] = 32'd2148021305;
        ram[69][127:96] = 32'd2094091315;
        ram[70][31:0] = 32'd1630538625;
        ram[70][63:32] = 32'd1777173702;
        ram[70][95:64] = 32'd618233280;
        ram[70][127:96] = 32'd3321912760;
        ram[71][31:0] = 32'd258676554;
        ram[71][63:32] = 32'd705180939;
        ram[71][95:64] = 32'd667168271;
        ram[71][127:96] = 32'd4136431290;
        ram[72][31:0] = 32'd262849900;
        ram[72][63:32] = 32'd496729428;
        ram[72][95:64] = 32'd3259086999;
        ram[72][127:96] = 32'd3072874000;
        ram[73][31:0] = 32'd3655331836;
        ram[73][63:32] = 32'd2329958859;
        ram[73][95:64] = 32'd2380132845;
        ram[73][127:96] = 32'd174084525;
        ram[74][31:0] = 32'd2975286243;
        ram[74][63:32] = 32'd141773217;
        ram[74][95:64] = 32'd265452422;
        ram[74][127:96] = 32'd3042141155;
        ram[75][31:0] = 32'd2360300364;
        ram[75][63:32] = 32'd3675695667;
        ram[75][95:64] = 32'd1076008577;
        ram[75][127:96] = 32'd3582560146;
        ram[76][31:0] = 32'd885943171;
        ram[76][63:32] = 32'd703237827;
        ram[76][95:64] = 32'd1771546382;
        ram[76][127:96] = 32'd66197177;
        ram[77][31:0] = 32'd1001871782;
        ram[77][63:32] = 32'd2815024490;
        ram[77][95:64] = 32'd4118581448;
        ram[77][127:96] = 32'd1351719823;
        ram[78][31:0] = 32'd1486852230;
        ram[78][63:32] = 32'd2976916899;
        ram[78][95:64] = 32'd4198757162;
        ram[78][127:96] = 32'd2804730422;
        ram[79][31:0] = 32'd1243284332;
        ram[79][63:32] = 32'd308852545;
        ram[79][95:64] = 32'd3083830815;
        ram[79][127:96] = 32'd2414245508;
        ram[80][31:0] = 32'd1627082053;
        ram[80][63:32] = 32'd3510587126;
        ram[80][95:64] = 32'd2713500914;
        ram[80][127:96] = 32'd650349116;
        ram[81][31:0] = 32'd3240530051;
        ram[81][63:32] = 32'd3825338226;
        ram[81][95:64] = 32'd626374968;
        ram[81][127:96] = 32'd614436650;
        ram[82][31:0] = 32'd1334801209;
        ram[82][63:32] = 32'd2440077942;
        ram[82][95:64] = 32'd2270922047;
        ram[82][127:96] = 32'd2402963099;
        ram[83][31:0] = 32'd3102777969;
        ram[83][63:32] = 32'd3264659335;
        ram[83][95:64] = 32'd4019955731;
        ram[83][127:96] = 32'd3512696420;
        ram[84][31:0] = 32'd2106753642;
        ram[84][63:32] = 32'd264400746;
        ram[84][95:64] = 32'd1698806919;
        ram[84][127:96] = 32'd3510710878;
        ram[85][31:0] = 32'd1961019814;
        ram[85][63:32] = 32'd720341552;
        ram[85][95:64] = 32'd1039652526;
        ram[85][127:96] = 32'd2034529216;
        ram[86][31:0] = 32'd2140186060;
        ram[86][63:32] = 32'd2552656500;
        ram[86][95:64] = 32'd1421834461;
        ram[86][127:96] = 32'd3262654288;
        ram[87][31:0] = 32'd2236840192;
        ram[87][63:32] = 32'd3136771072;
        ram[87][95:64] = 32'd3916124113;
        ram[87][127:96] = 32'd4052137824;
        ram[88][31:0] = 32'd1475447480;
        ram[88][63:32] = 32'd1320710077;
        ram[88][95:64] = 32'd1554725479;
        ram[88][127:96] = 32'd2340500150;
        ram[89][31:0] = 32'd2499526742;
        ram[89][63:32] = 32'd2986504088;
        ram[89][95:64] = 32'd3518005260;
        ram[89][127:96] = 32'd3381025996;
        ram[90][31:0] = 32'd3720302651;
        ram[90][63:32] = 32'd3093348283;
        ram[90][95:64] = 32'd1169309859;
        ram[90][127:96] = 32'd3448701357;
        ram[91][31:0] = 32'd3098727765;
        ram[91][63:32] = 32'd4037880385;
        ram[91][95:64] = 32'd2558372418;
        ram[91][127:96] = 32'd3102588231;
        ram[92][31:0] = 32'd329657286;
        ram[92][63:32] = 32'd3108046467;
        ram[92][95:64] = 32'd4079085858;
        ram[92][127:96] = 32'd2128993578;
        ram[93][31:0] = 32'd1694808878;
        ram[93][63:32] = 32'd843400262;
        ram[93][95:64] = 32'd3344969860;
        ram[93][127:96] = 32'd116681397;
        ram[94][31:0] = 32'd2751670357;
        ram[94][63:32] = 32'd385500254;
        ram[94][95:64] = 32'd1591577112;
        ram[94][127:96] = 32'd3734682012;
        ram[95][31:0] = 32'd3066489922;
        ram[95][63:32] = 32'd3015459872;
        ram[95][95:64] = 32'd3756847522;
        ram[95][127:96] = 32'd1615749578;
        ram[96][31:0] = 32'd2950368077;
        ram[96][63:32] = 32'd362704286;
        ram[96][95:64] = 32'd1528358932;
        ram[96][127:96] = 32'd2723287972;
        ram[97][31:0] = 32'd1640297598;
        ram[97][63:32] = 32'd4254260300;
        ram[97][95:64] = 32'd1994867427;
        ram[97][127:96] = 32'd3059314876;
        ram[98][31:0] = 32'd1235012268;
        ram[98][63:32] = 32'd3328956941;
        ram[98][95:64] = 32'd438437706;
        ram[98][127:96] = 32'd1385063468;
        ram[99][31:0] = 32'd2144452371;
        ram[99][63:32] = 32'd1685622093;
        ram[99][95:64] = 32'd31940929;
        ram[99][127:96] = 32'd2238490792;
        ram[100][31:0] = 32'd361266538;
        ram[100][63:32] = 32'd1922832907;
        ram[100][95:64] = 32'd4154520894;
        ram[100][127:96] = 32'd1005991444;
        ram[101][31:0] = 32'd586528649;
        ram[101][63:32] = 32'd3625043014;
        ram[101][95:64] = 32'd3304677203;
        ram[101][127:96] = 32'd1151535682;
        ram[102][31:0] = 32'd303432423;
        ram[102][63:32] = 32'd1379904639;
        ram[102][95:64] = 32'd3327850702;
        ram[102][127:96] = 32'd3771831217;
        ram[103][31:0] = 32'd38261169;
        ram[103][63:32] = 32'd4153973033;
        ram[103][95:64] = 32'd998493570;
        ram[103][127:96] = 32'd1573085486;
        ram[104][31:0] = 32'd593392457;
        ram[104][63:32] = 32'd2340832447;
        ram[104][95:64] = 32'd1103181938;
        ram[104][127:96] = 32'd2926357254;
        ram[105][31:0] = 32'd3361591300;
        ram[105][63:32] = 32'd3457007363;
        ram[105][95:64] = 32'd533866239;
        ram[105][127:96] = 32'd3386031789;
        ram[106][31:0] = 32'd1637986519;
        ram[106][63:32] = 32'd3413574269;
        ram[106][95:64] = 32'd1898868723;
        ram[106][127:96] = 32'd3283430231;
        ram[107][31:0] = 32'd5484622;
        ram[107][63:32] = 32'd1861495304;
        ram[107][95:64] = 32'd863164190;
        ram[107][127:96] = 32'd1733952639;
        ram[108][31:0] = 32'd3643494175;
        ram[108][63:32] = 32'd764669096;
        ram[108][95:64] = 32'd425295928;
        ram[108][127:96] = 32'd2086475014;
        ram[109][31:0] = 32'd3704035340;
        ram[109][63:32] = 32'd2756765652;
        ram[109][95:64] = 32'd3272117358;
        ram[109][127:96] = 32'd3398516884;
        ram[110][31:0] = 32'd1696256247;
        ram[110][63:32] = 32'd948216216;
        ram[110][95:64] = 32'd659523681;
        ram[110][127:96] = 32'd3697129869;
        ram[111][31:0] = 32'd2818036757;
        ram[111][63:32] = 32'd495816375;
        ram[111][95:64] = 32'd1055605986;
        ram[111][127:96] = 32'd1438660782;
        ram[112][31:0] = 32'd738342312;
        ram[112][63:32] = 32'd3226103403;
        ram[112][95:64] = 32'd2465959336;
        ram[112][127:96] = 32'd903750376;
        ram[113][31:0] = 32'd4242215536;
        ram[113][63:32] = 32'd3500901833;
        ram[113][95:64] = 32'd885130039;
        ram[113][127:96] = 32'd442340444;
        ram[114][31:0] = 32'd2194731325;
        ram[114][63:32] = 32'd4191839408;
        ram[114][95:64] = 32'd4229334037;
        ram[114][127:96] = 32'd1569664529;
        ram[115][31:0] = 32'd544566434;
        ram[115][63:32] = 32'd2300259007;
        ram[115][95:64] = 32'd1029956024;
        ram[115][127:96] = 32'd358187220;
        ram[116][31:0] = 32'd1513902136;
        ram[116][63:32] = 32'd4289052588;
        ram[116][95:64] = 32'd3439948819;
        ram[116][127:96] = 32'd3833684444;
        ram[117][31:0] = 32'd631997243;
        ram[117][63:32] = 32'd421173559;
        ram[117][95:64] = 32'd4198953116;
        ram[117][127:96] = 32'd3963935252;
        ram[118][31:0] = 32'd3690519590;
        ram[118][63:32] = 32'd893693086;
        ram[118][95:64] = 32'd3709210581;
        ram[118][127:96] = 32'd1268256802;
        ram[119][31:0] = 32'd1210849249;
        ram[119][63:32] = 32'd2712954145;
        ram[119][95:64] = 32'd2214102913;
        ram[119][127:96] = 32'd3387098527;
        ram[120][31:0] = 32'd2118543923;
        ram[120][63:32] = 32'd1841367641;
        ram[120][95:64] = 32'd931171768;
        ram[120][127:96] = 32'd1127608633;
        ram[121][31:0] = 32'd3316009856;
        ram[121][63:32] = 32'd4058835011;
        ram[121][95:64] = 32'd3076352410;
        ram[121][127:96] = 32'd1196914595;
        ram[122][31:0] = 32'd3891522968;
        ram[122][63:32] = 32'd4219814471;
        ram[122][95:64] = 32'd309980754;
        ram[122][127:96] = 32'd1350952293;
        ram[123][31:0] = 32'd3279720460;
        ram[123][63:32] = 32'd2901124810;
        ram[123][95:64] = 32'd1860698751;
        ram[123][127:96] = 32'd2224122238;
        ram[124][31:0] = 32'd2547440168;
        ram[124][63:32] = 32'd2929216944;
        ram[124][95:64] = 32'd1844922442;
        ram[124][127:96] = 32'd3027405431;
        ram[125][31:0] = 32'd1137385221;
        ram[125][63:32] = 32'd138578467;
        ram[125][95:64] = 32'd1213399919;
        ram[125][127:96] = 32'd3936231662;
        ram[126][31:0] = 32'd3287718623;
        ram[126][63:32] = 32'd3673032087;
        ram[126][95:64] = 32'd659028168;
        ram[126][127:96] = 32'd3886571279;
        ram[127][31:0] = 32'd2458412144;
        ram[127][63:32] = 32'd2005844869;
        ram[127][95:64] = 32'd195368792;
        ram[127][127:96] = 32'd3832262737;
        ram[128][31:0] = 32'd3640518258;
        ram[128][63:32] = 32'd2469969087;
        ram[128][95:64] = 32'd1369178089;
        ram[128][127:96] = 32'd810273649;
        ram[129][31:0] = 32'd3801022005;
        ram[129][63:32] = 32'd301926624;
        ram[129][95:64] = 32'd4044851709;
        ram[129][127:96] = 32'd818470911;
        ram[130][31:0] = 32'd2738263273;
        ram[130][63:32] = 32'd251937582;
        ram[130][95:64] = 32'd160969124;
        ram[130][127:96] = 32'd662160688;
        ram[131][31:0] = 32'd527412138;
        ram[131][63:32] = 32'd2405063111;
        ram[131][95:64] = 32'd512884825;
        ram[131][127:96] = 32'd3071282313;
        ram[132][31:0] = 32'd779927443;
        ram[132][63:32] = 32'd3797362521;
        ram[132][95:64] = 32'd3894234752;
        ram[132][127:96] = 32'd1030173785;
        ram[133][31:0] = 32'd720228296;
        ram[133][63:32] = 32'd79829296;
        ram[133][95:64] = 32'd909548475;
        ram[133][127:96] = 32'd3322326490;
        ram[134][31:0] = 32'd1287154060;
        ram[134][63:32] = 32'd1818603648;
        ram[134][95:64] = 32'd3291868179;
        ram[134][127:96] = 32'd2220181209;
        ram[135][31:0] = 32'd3411388360;
        ram[135][63:32] = 32'd2903716974;
        ram[135][95:64] = 32'd1293852496;
        ram[135][127:96] = 32'd1828813246;
        ram[136][31:0] = 32'd3425081071;
        ram[136][63:32] = 32'd2528965743;
        ram[136][95:64] = 32'd3391432801;
        ram[136][127:96] = 32'd2078655512;
        ram[137][31:0] = 32'd1224644377;
        ram[137][63:32] = 32'd3183535881;
        ram[137][95:64] = 32'd4137090125;
        ram[137][127:96] = 32'd2595070212;
        ram[138][31:0] = 32'd1826755672;
        ram[138][63:32] = 32'd255303072;
        ram[138][95:64] = 32'd2441644451;
        ram[138][127:96] = 32'd656657158;
        ram[139][31:0] = 32'd1863958673;
        ram[139][63:32] = 32'd584829879;
        ram[139][95:64] = 32'd1054185022;
        ram[139][127:96] = 32'd4164214068;
        ram[140][31:0] = 32'd2283876130;
        ram[140][63:32] = 32'd1153481128;
        ram[140][95:64] = 32'd3051066239;
        ram[140][127:96] = 32'd3249157073;
        ram[141][31:0] = 32'd1053780301;
        ram[141][63:32] = 32'd3726381274;
        ram[141][95:64] = 32'd3343708057;
        ram[141][127:96] = 32'd1569593133;
        ram[142][31:0] = 32'd3549289617;
        ram[142][63:32] = 32'd2945905132;
        ram[142][95:64] = 32'd1605140899;
        ram[142][127:96] = 32'd2093197089;
        ram[143][31:0] = 32'd2425967003;
        ram[143][63:32] = 32'd3896166626;
        ram[143][95:64] = 32'd164286464;
        ram[143][127:96] = 32'd2983705835;
        ram[144][31:0] = 32'd3615860568;
        ram[144][63:32] = 32'd2874325634;
        ram[144][95:64] = 32'd7656595;
        ram[144][127:96] = 32'd2251069002;
        ram[145][31:0] = 32'd4090953264;
        ram[145][63:32] = 32'd1862601448;
        ram[145][95:64] = 32'd3203865679;
        ram[145][127:96] = 32'd2629654119;
        ram[146][31:0] = 32'd488666373;
        ram[146][63:32] = 32'd3271570656;
        ram[146][95:64] = 32'd441018196;
        ram[146][127:96] = 32'd398702022;
        ram[147][31:0] = 32'd2588161959;
        ram[147][63:32] = 32'd150013310;
        ram[147][95:64] = 32'd4086930734;
        ram[147][127:96] = 32'd2185077938;
        ram[148][31:0] = 32'd531026440;
        ram[148][63:32] = 32'd4289367533;
        ram[148][95:64] = 32'd3713092353;
        ram[148][127:96] = 32'd2353985372;
        ram[149][31:0] = 32'd1619445656;
        ram[149][63:32] = 32'd2521741564;
        ram[149][95:64] = 32'd402461654;
        ram[149][127:96] = 32'd2679728859;
        ram[150][31:0] = 32'd2274691543;
        ram[150][63:32] = 32'd1792044048;
        ram[150][95:64] = 32'd3974529998;
        ram[150][127:96] = 32'd631643568;
        ram[151][31:0] = 32'd1821330664;
        ram[151][63:32] = 32'd3854904784;
        ram[151][95:64] = 32'd1654540681;
        ram[151][127:96] = 32'd2212965614;
        ram[152][31:0] = 32'd3588334251;
        ram[152][63:32] = 32'd779641857;
        ram[152][95:64] = 32'd4072126458;
        ram[152][127:96] = 32'd1073177235;
        ram[153][31:0] = 32'd1343092192;
        ram[153][63:32] = 32'd1975594517;
        ram[153][95:64] = 32'd292281791;
        ram[153][127:96] = 32'd3415332789;
        ram[154][31:0] = 32'd1933938369;
        ram[154][63:32] = 32'd306081816;
        ram[154][95:64] = 32'd2836784331;
        ram[154][127:96] = 32'd3534431847;
        ram[155][31:0] = 32'd990877164;
        ram[155][63:32] = 32'd2700116951;
        ram[155][95:64] = 32'd981558266;
        ram[155][127:96] = 32'd1100459140;
        ram[156][31:0] = 32'd3685889770;
        ram[156][63:32] = 32'd402550184;
        ram[156][95:64] = 32'd1133261423;
        ram[156][127:96] = 32'd2656035837;
        ram[157][31:0] = 32'd2527456798;
        ram[157][63:32] = 32'd701803144;
        ram[157][95:64] = 32'd1885255059;
        ram[157][127:96] = 32'd1893022681;
        ram[158][31:0] = 32'd1155677548;
        ram[158][63:32] = 32'd1648345772;
        ram[158][95:64] = 32'd829790260;
        ram[158][127:96] = 32'd2467999083;
        ram[159][31:0] = 32'd1043611674;
        ram[159][63:32] = 32'd2030896509;
        ram[159][95:64] = 32'd2536119541;
        ram[159][127:96] = 32'd3943965978;
        ram[160][31:0] = 32'd2917644381;
        ram[160][63:32] = 32'd2076475850;
        ram[160][95:64] = 32'd2479303443;
        ram[160][127:96] = 32'd4288523406;
        ram[161][31:0] = 32'd2060679594;
        ram[161][63:32] = 32'd1184230149;
        ram[161][95:64] = 32'd132734761;
        ram[161][127:96] = 32'd1466466644;
        ram[162][31:0] = 32'd2126227131;
        ram[162][63:32] = 32'd3331514741;
        ram[162][95:64] = 32'd621028655;
        ram[162][127:96] = 32'd1407051673;
        ram[163][31:0] = 32'd3031069961;
        ram[163][63:32] = 32'd2828538946;
        ram[163][95:64] = 32'd3194778842;
        ram[163][127:96] = 32'd300940477;
        ram[164][31:0] = 32'd2417503440;
        ram[164][63:32] = 32'd927834072;
        ram[164][95:64] = 32'd2510800920;
        ram[164][127:96] = 32'd3342857150;
        ram[165][31:0] = 32'd2333695448;
        ram[165][63:32] = 32'd2978772408;
        ram[165][95:64] = 32'd2797788974;
        ram[165][127:96] = 32'd367404024;
        ram[166][31:0] = 32'd836176777;
        ram[166][63:32] = 32'd864347332;
        ram[166][95:64] = 32'd788353255;
        ram[166][127:96] = 32'd3439559431;
        ram[167][31:0] = 32'd1703734548;
        ram[167][63:32] = 32'd459165770;
        ram[167][95:64] = 32'd5269375;
        ram[167][127:96] = 32'd3933977752;
        ram[168][31:0] = 32'd1691338492;
        ram[168][63:32] = 32'd102644394;
        ram[168][95:64] = 32'd1833629200;
        ram[168][127:96] = 32'd2346375170;
        ram[169][31:0] = 32'd1600125893;
        ram[169][63:32] = 32'd73624117;
        ram[169][95:64] = 32'd3688685586;
        ram[169][127:96] = 32'd2092664236;
        ram[170][31:0] = 32'd555640076;
        ram[170][63:32] = 32'd2735001250;
        ram[170][95:64] = 32'd3207157459;
        ram[170][127:96] = 32'd3125603621;
        ram[171][31:0] = 32'd4096736423;
        ram[171][63:32] = 32'd2966388477;
        ram[171][95:64] = 32'd4286094390;
        ram[171][127:96] = 32'd1851326025;
        ram[172][31:0] = 32'd3601440211;
        ram[172][63:32] = 32'd753035072;
        ram[172][95:64] = 32'd4288616562;
        ram[172][127:96] = 32'd3704402127;
        ram[173][31:0] = 32'd142573271;
        ram[173][63:32] = 32'd107943679;
        ram[173][95:64] = 32'd11288168;
        ram[173][127:96] = 32'd650862610;
        ram[174][31:0] = 32'd3092369021;
        ram[174][63:32] = 32'd1149613355;
        ram[174][95:64] = 32'd3118469034;
        ram[174][127:96] = 32'd1874804212;
        ram[175][31:0] = 32'd2118661662;
        ram[175][63:32] = 32'd202904808;
        ram[175][95:64] = 32'd2449747273;
        ram[175][127:96] = 32'd3644357459;
        ram[176][31:0] = 32'd2828619334;
        ram[176][63:32] = 32'd3595301892;
        ram[176][95:64] = 32'd2740353206;
        ram[176][127:96] = 32'd1855980571;
        ram[177][31:0] = 32'd4183077687;
        ram[177][63:32] = 32'd2882321478;
        ram[177][95:64] = 32'd2873504019;
        ram[177][127:96] = 32'd2188493423;
        ram[178][31:0] = 32'd3498676098;
        ram[178][63:32] = 32'd358436771;
        ram[178][95:64] = 32'd4030058467;
        ram[178][127:96] = 32'd662596021;
        ram[179][31:0] = 32'd2231466293;
        ram[179][63:32] = 32'd3753177976;
        ram[179][95:64] = 32'd471550192;
        ram[179][127:96] = 32'd1608144627;
        ram[180][31:0] = 32'd3049260861;
        ram[180][63:32] = 32'd3714234635;
        ram[180][95:64] = 32'd3788823028;
        ram[180][127:96] = 32'd2519917846;
        ram[181][31:0] = 32'd2951008079;
        ram[181][63:32] = 32'd383602951;
        ram[181][95:64] = 32'd750377268;
        ram[181][127:96] = 32'd2548078876;
        ram[182][31:0] = 32'd820874592;
        ram[182][63:32] = 32'd1893345796;
        ram[182][95:64] = 32'd237210761;
        ram[182][127:96] = 32'd4083566603;
        ram[183][31:0] = 32'd1612454682;
        ram[183][63:32] = 32'd1395512612;
        ram[183][95:64] = 32'd2662220977;
        ram[183][127:96] = 32'd662603260;
        ram[184][31:0] = 32'd4060815809;
        ram[184][63:32] = 32'd1797063890;
        ram[184][95:64] = 32'd2491419620;
        ram[184][127:96] = 32'd24113143;
        ram[185][31:0] = 32'd3140061557;
        ram[185][63:32] = 32'd1930615449;
        ram[185][95:64] = 32'd3025146857;
        ram[185][127:96] = 32'd1004600950;
        ram[186][31:0] = 32'd2105270382;
        ram[186][63:32] = 32'd2968700236;
        ram[186][95:64] = 32'd1047595471;
        ram[186][127:96] = 32'd3403950629;
        ram[187][31:0] = 32'd2905536779;
        ram[187][63:32] = 32'd1442235455;
        ram[187][95:64] = 32'd86667935;
        ram[187][127:96] = 32'd616267458;
        ram[188][31:0] = 32'd2638568597;
        ram[188][63:32] = 32'd3408944389;
        ram[188][95:64] = 32'd2262784563;
        ram[188][127:96] = 32'd1863651176;
        ram[189][31:0] = 32'd701769280;
        ram[189][63:32] = 32'd1051045639;
        ram[189][95:64] = 32'd2116480522;
        ram[189][127:96] = 32'd2171230616;
        ram[190][31:0] = 32'd1471651428;
        ram[190][63:32] = 32'd1203634462;
        ram[190][95:64] = 32'd2385791137;
        ram[190][127:96] = 32'd1119246121;
        ram[191][31:0] = 32'd3790187111;
        ram[191][63:32] = 32'd3971243364;
        ram[191][95:64] = 32'd3995767260;
        ram[191][127:96] = 32'd1189601977;
        ram[192][31:0] = 32'd499123626;
        ram[192][63:32] = 32'd1388272500;
        ram[192][95:64] = 32'd2171678767;
        ram[192][127:96] = 32'd733190410;
        ram[193][31:0] = 32'd925346153;
        ram[193][63:32] = 32'd531933772;
        ram[193][95:64] = 32'd2834186409;
        ram[193][127:96] = 32'd1482893985;
        ram[194][31:0] = 32'd1107570546;
        ram[194][63:32] = 32'd850545293;
        ram[194][95:64] = 32'd75381009;
        ram[194][127:96] = 32'd1944019024;
        ram[195][31:0] = 32'd614300779;
        ram[195][63:32] = 32'd1625107923;
        ram[195][95:64] = 32'd3267113827;
        ram[195][127:96] = 32'd1379073191;
        ram[196][31:0] = 32'd1428448895;
        ram[196][63:32] = 32'd1809300641;
        ram[196][95:64] = 32'd3135983681;
        ram[196][127:96] = 32'd2332338642;
        ram[197][31:0] = 32'd3488647823;
        ram[197][63:32] = 32'd1966886339;
        ram[197][95:64] = 32'd3349018487;
        ram[197][127:96] = 32'd1872473622;
        ram[198][31:0] = 32'd758407755;
        ram[198][63:32] = 32'd3367465369;
        ram[198][95:64] = 32'd1845668888;
        ram[198][127:96] = 32'd88944858;
        ram[199][31:0] = 32'd1296508384;
        ram[199][63:32] = 32'd3094034019;
        ram[199][95:64] = 32'd606531690;
        ram[199][127:96] = 32'd3141851948;
        ram[200][31:0] = 32'd3860457312;
        ram[200][63:32] = 32'd991402029;
        ram[200][95:64] = 32'd3968035631;
        ram[200][127:96] = 32'd3117956401;
        ram[201][31:0] = 32'd493963406;
        ram[201][63:32] = 32'd2845628761;
        ram[201][95:64] = 32'd581402204;
        ram[201][127:96] = 32'd381283231;
        ram[202][31:0] = 32'd4052309515;
        ram[202][63:32] = 32'd3862961053;
        ram[202][95:64] = 32'd1470816688;
        ram[202][127:96] = 32'd3068252576;
        ram[203][31:0] = 32'd2158247624;
        ram[203][63:32] = 32'd2639132952;
        ram[203][95:64] = 32'd3975966587;
        ram[203][127:96] = 32'd2868329003;
        ram[204][31:0] = 32'd2846493614;
        ram[204][63:32] = 32'd3133004597;
        ram[204][95:64] = 32'd3235329560;
        ram[204][127:96] = 32'd1751705146;
        ram[205][31:0] = 32'd2100567583;
        ram[205][63:32] = 32'd4085841762;
        ram[205][95:64] = 32'd2970417653;
        ram[205][127:96] = 32'd700710660;
        ram[206][31:0] = 32'd403117584;
        ram[206][63:32] = 32'd4252998212;
        ram[206][95:64] = 32'd4190783551;
        ram[206][127:96] = 32'd1675509145;
        ram[207][31:0] = 32'd3426927664;
        ram[207][63:32] = 32'd1714014072;
        ram[207][95:64] = 32'd639045237;
        ram[207][127:96] = 32'd3525708661;
        ram[208][31:0] = 32'd1247309753;
        ram[208][63:32] = 32'd2181837440;
        ram[208][95:64] = 32'd2481571039;
        ram[208][127:96] = 32'd4032415179;
        ram[209][31:0] = 32'd2452486217;
        ram[209][63:32] = 32'd1693487156;
        ram[209][95:64] = 32'd4110932613;
        ram[209][127:96] = 32'd1534108225;
        ram[210][31:0] = 32'd2554070727;
        ram[210][63:32] = 32'd1919489441;
        ram[210][95:64] = 32'd4112986047;
        ram[210][127:96] = 32'd1944986852;
        ram[211][31:0] = 32'd883501816;
        ram[211][63:32] = 32'd4092281317;
        ram[211][95:64] = 32'd2824502397;
        ram[211][127:96] = 32'd1925753163;
        ram[212][31:0] = 32'd74868948;
        ram[212][63:32] = 32'd2242143770;
        ram[212][95:64] = 32'd2610616633;
        ram[212][127:96] = 32'd1149027704;
        ram[213][31:0] = 32'd443188871;
        ram[213][63:32] = 32'd3949017632;
        ram[213][95:64] = 32'd2209713226;
        ram[213][127:96] = 32'd2722662011;
        ram[214][31:0] = 32'd4086119564;
        ram[214][63:32] = 32'd1114468449;
        ram[214][95:64] = 32'd1864704728;
        ram[214][127:96] = 32'd951891562;
        ram[215][31:0] = 32'd4017842051;
        ram[215][63:32] = 32'd3560847281;
        ram[215][95:64] = 32'd1375551832;
        ram[215][127:96] = 32'd1442050635;
        ram[216][31:0] = 32'd702666674;
        ram[216][63:32] = 32'd2216532256;
        ram[216][95:64] = 32'd2280351118;
        ram[216][127:96] = 32'd3206650022;
        ram[217][31:0] = 32'd2145195459;
        ram[217][63:32] = 32'd707255610;
        ram[217][95:64] = 32'd939174474;
        ram[217][127:96] = 32'd1185961275;
        ram[218][31:0] = 32'd1431148747;
        ram[218][63:32] = 32'd1792266633;
        ram[218][95:64] = 32'd3881945575;
        ram[218][127:96] = 32'd717937086;
        ram[219][31:0] = 32'd3195243728;
        ram[219][63:32] = 32'd4061042516;
        ram[219][95:64] = 32'd1635543175;
        ram[219][127:96] = 32'd978943048;
        ram[220][31:0] = 32'd1460846078;
        ram[220][63:32] = 32'd3445283547;
        ram[220][95:64] = 32'd1957393229;
        ram[220][127:96] = 32'd43240007;
        ram[221][31:0] = 32'd678817658;
        ram[221][63:32] = 32'd1024871351;
        ram[221][95:64] = 32'd479387173;
        ram[221][127:96] = 32'd852431783;
        ram[222][31:0] = 32'd2075271081;
        ram[222][63:32] = 32'd3384816046;
        ram[222][95:64] = 32'd1732209976;
        ram[222][127:96] = 32'd2459813267;
        ram[223][31:0] = 32'd2706547949;
        ram[223][63:32] = 32'd3704026762;
        ram[223][95:64] = 32'd844419571;
        ram[223][127:96] = 32'd2712734655;
        ram[224][31:0] = 32'd3066857618;
        ram[224][63:32] = 32'd1039575909;
        ram[224][95:64] = 32'd3668671927;
        ram[224][127:96] = 32'd2738438795;
        ram[225][31:0] = 32'd2793424475;
        ram[225][63:32] = 32'd2235022597;
        ram[225][95:64] = 32'd378352142;
        ram[225][127:96] = 32'd3268229861;
        ram[226][31:0] = 32'd4135674155;
        ram[226][63:32] = 32'd444182793;
        ram[226][95:64] = 32'd3294149566;
        ram[226][127:96] = 32'd2677761354;
        ram[227][31:0] = 32'd192450639;
        ram[227][63:32] = 32'd1277973101;
        ram[227][95:64] = 32'd3948715188;
        ram[227][127:96] = 32'd949505153;
        ram[228][31:0] = 32'd1730083639;
        ram[228][63:32] = 32'd81643281;
        ram[228][95:64] = 32'd336515192;
        ram[228][127:96] = 32'd275549499;
        ram[229][31:0] = 32'd379022188;
        ram[229][63:32] = 32'd778607413;
        ram[229][95:64] = 32'd3205683197;
        ram[229][127:96] = 32'd4037234632;
        ram[230][31:0] = 32'd1092104427;
        ram[230][63:32] = 32'd2725134890;
        ram[230][95:64] = 32'd3546517031;
        ram[230][127:96] = 32'd412824823;
        ram[231][31:0] = 32'd2722183945;
        ram[231][63:32] = 32'd1219013972;
        ram[231][95:64] = 32'd2655641510;
        ram[231][127:96] = 32'd1780961405;
        ram[232][31:0] = 32'd3416090981;
        ram[232][63:32] = 32'd2524469636;
        ram[232][95:64] = 32'd528430591;
        ram[232][127:96] = 32'd12882843;
        ram[233][31:0] = 32'd1138021835;
        ram[233][63:32] = 32'd1333871334;
        ram[233][95:64] = 32'd3429994139;
        ram[233][127:96] = 32'd1724373865;
        ram[234][31:0] = 32'd1292504590;
        ram[234][63:32] = 32'd1789369773;
        ram[234][95:64] = 32'd2569444219;
        ram[234][127:96] = 32'd3724952086;
        ram[235][31:0] = 32'd1592502160;
        ram[235][63:32] = 32'd4153701105;
        ram[235][95:64] = 32'd916379260;
        ram[235][127:96] = 32'd2355932002;
        ram[236][31:0] = 32'd2878291750;
        ram[236][63:32] = 32'd3470321335;
        ram[236][95:64] = 32'd88830842;
        ram[236][127:96] = 32'd3401316327;
        ram[237][31:0] = 32'd2974746974;
        ram[237][63:32] = 32'd1115900148;
        ram[237][95:64] = 32'd1338640197;
        ram[237][127:96] = 32'd2460043506;
        ram[238][31:0] = 32'd4122296222;
        ram[238][63:32] = 32'd1006062678;
        ram[238][95:64] = 32'd643086006;
        ram[238][127:96] = 32'd1186627500;
        ram[239][31:0] = 32'd2021668976;
        ram[239][63:32] = 32'd1537653831;
        ram[239][95:64] = 32'd1861866575;
        ram[239][127:96] = 32'd88139643;
        ram[240][31:0] = 32'd2916006627;
        ram[240][63:32] = 32'd1106788918;
        ram[240][95:64] = 32'd1878395484;
        ram[240][127:96] = 32'd11250872;
        ram[241][31:0] = 32'd3846880485;
        ram[241][63:32] = 32'd2839272030;
        ram[241][95:64] = 32'd4123438644;
        ram[241][127:96] = 32'd4013713639;
        ram[242][31:0] = 32'd2279943055;
        ram[242][63:32] = 32'd211093134;
        ram[242][95:64] = 32'd3921400631;
        ram[242][127:96] = 32'd1742952547;
        ram[243][31:0] = 32'd2852470675;
        ram[243][63:32] = 32'd251047168;
        ram[243][95:64] = 32'd4232010606;
        ram[243][127:96] = 32'd3780880889;
        ram[244][31:0] = 32'd1630561231;
        ram[244][63:32] = 32'd4221183128;
        ram[244][95:64] = 32'd1849704765;
        ram[244][127:96] = 32'd1293811238;
        ram[245][31:0] = 32'd951388280;
        ram[245][63:32] = 32'd1037042201;
        ram[245][95:64] = 32'd441351460;
        ram[245][127:96] = 32'd3867328918;
        ram[246][31:0] = 32'd2904690682;
        ram[246][63:32] = 32'd212834635;
        ram[246][95:64] = 32'd942798349;
        ram[246][127:96] = 32'd4200030814;
        ram[247][31:0] = 32'd2921234412;
        ram[247][63:32] = 32'd2993705083;
        ram[247][95:64] = 32'd616895957;
        ram[247][127:96] = 32'd1186657120;
        ram[248][31:0] = 32'd660776973;
        ram[248][63:32] = 32'd2081880215;
        ram[248][95:64] = 32'd2394012061;
        ram[248][127:96] = 32'd2930137711;
        ram[249][31:0] = 32'd3896560801;
        ram[249][63:32] = 32'd2373012430;
        ram[249][95:64] = 32'd4165651510;
        ram[249][127:96] = 32'd3554282325;
        ram[250][31:0] = 32'd3122678110;
        ram[250][63:32] = 32'd2446236361;
        ram[250][95:64] = 32'd800960759;
        ram[250][127:96] = 32'd3015381937;
        ram[251][31:0] = 32'd2043377402;
        ram[251][63:32] = 32'd3281370832;
        ram[251][95:64] = 32'd1278342728;
        ram[251][127:96] = 32'd240134872;
        ram[252][31:0] = 32'd3635208870;
        ram[252][63:32] = 32'd1069602971;
        ram[252][95:64] = 32'd70305260;
        ram[252][127:96] = 32'd3132942458;
        ram[253][31:0] = 32'd3611161271;
        ram[253][63:32] = 32'd3443847325;
        ram[253][95:64] = 32'd2402115690;
        ram[253][127:96] = 32'd2967419399;
        ram[254][31:0] = 32'd1576676339;
        ram[254][63:32] = 32'd770943859;
        ram[254][95:64] = 32'd1157429103;
        ram[254][127:96] = 32'd510091675;
        ram[255][31:0] = 32'd3144327154;
        ram[255][63:32] = 32'd2654480329;
        ram[255][95:64] = 32'd3690728159;
        ram[255][127:96] = 32'd107160650;

    end
    always @(posedge clk) begin
        addr_r <= raddr;
        if(we) ram[waddr] <= din;
    end
    assign dout = ram[addr_r]; 

endmodule
