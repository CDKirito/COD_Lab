
/*
本文件是一个测试文件，用于测试cache模块
工作原理是模仿CPU的读写请求，对cache进行读写操作
将Cache返回的数据与预先数据进行比较，如果一致则测试通过
*/
`timescale 1ns/1ps
module cache_tb();

    //测试参数
    parameter READ_NUM = 2000;  // 测试次数 这里设置为2000次读，1000次写
    parameter WRITE_NUM = 1000;  
    //模块参数
    parameter INDEX_WIDTH       = 3;   // Cache索引位宽 2^3=8行
    parameter LINE_OFFSET_WIDTH = 2;   // 行偏移位宽，决定了一行的宽度 2^2=4字
    parameter SPACE_OFFSET      = 2;   // 一个地址空间占1个字节，因此一个字需要4个地址空间，由于假设为整字读取，处理地址的时候可以默认后两位为0
    parameter MEM_ADDR_WIDTH    = 10;   // 为了简化，这里假设内存地址宽度为10位（CPU请求地址仍然是32位，只不过我们这里简化处理，截断了高位） 
    parameter WAY_NUM           = 4;   // Cache N路组相联(N=1的时候是直接映射)

    // 变化的信号 CPU发出
    reg clk=1;
    reg rstn=1;
    reg stat=0;
    // 等rstn信号稳定后 clk信号才开始翻转
    initial begin
        #1 rstn = 0;
        #1 rstn = 1;
        stat = 1;
    end
    always  #1 clk = ~clk;

    wire [31:0] addr;
    wire r_req;
    wire w_req;
    wire [31:0] w_data;

    // 导线
    wire [31:0] r_data;
    wire miss;
    wire mem_r;
    wire mem_w;
    wire [31:0] mem_addr;
    wire [127:0] mem_w_data;
    wire [127:0] mem_r_data;
    wire mem_ready;

    // 用于测试的信号
    reg [MEM_ADDR_WIDTH-1:0] test_addr[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试地址
    reg [32:0] test_data[0:READ_NUM+WRITE_NUM-1];  // 用于存储测试数据 最高位用于标记是否写入 0：读 1：写
    reg [31:0] test_cnt=0;  // 用于计数，每次读写操作后加1
    reg diff=0;  // 用于标记是否有不一致的数据

    // 用于对比的提交，当前cache应该给出的数据
    wire op;
    wire[31:0] data;
    assign op = test_data[test_cnt-1][32];
    assign data = test_data[test_cnt-1][31:0];
    
    // 状态机
    assign addr = test_addr[test_cnt]<<SPACE_OFFSET;
    assign r_req = test_data[test_cnt][32] == 0 ? 1 : 0;
    assign w_req = test_data[test_cnt][32] == 1 ? 1 : 0;
    assign w_data = test_data[test_cnt][31:0];
    always @(posedge clk) begin
        if (!miss && (test_cnt < READ_NUM+WRITE_NUM) && stat) begin
            if (test_data[test_cnt-1][32] == 0) begin  // 读
                if (r_data != test_data[test_cnt-1][31:0]) begin
                    $display("Read error at %d, expect %h, get %h", test_cnt, test_data[test_cnt-1][31:0], r_data);
                    diff = 1;
                end
            end
            test_cnt <= test_cnt + 1;
        end
    end

    // 例化cache
    cache #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .WAY_NUM(WAY_NUM)
    ) cache_inst(
        .clk(clk),
        .rstn(rstn),
        .addr(addr),
        .r_req(r_req),
        .w_req(w_req),
        .w_data(w_data),
        .r_data(r_data),
        .miss(miss),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 内存
    mem #(
        .INDEX_WIDTH(INDEX_WIDTH),
        .LINE_OFFSET_WIDTH(LINE_OFFSET_WIDTH),
        .SPACE_OFFSET(SPACE_OFFSET),
        .MEM_ADDR_WIDTH(MEM_ADDR_WIDTH-LINE_OFFSET_WIDTH),
        .WAY_NUM(WAY_NUM)
    ) mem_inst(
        .clk(clk),
        .rstn(rstn),
        .mem_r(mem_r),
        .mem_w(mem_w),
        .mem_addr(mem_addr),
        .mem_w_data(mem_w_data),
        .mem_r_data(mem_r_data),
        .mem_ready(mem_ready)
    );

    // 初始化测试数据
    initial begin
        test_addr[0] = 907;
        test_data[0] = 33'd2677761354;
        test_addr[1] = 730;
        test_data[1] = 33'd237210761;
        test_addr[2] = 662;
        test_data[2] = 33'd7491117030;
        test_addr[3] = 666;
        test_data[3] = 33'd5743769147;
        test_addr[4] = 202;
        test_data[4] = 33'd3541495957;
        test_addr[5] = 271;
        test_data[5] = 33'd3753349860;
        test_addr[6] = 143;
        test_data[6] = 33'd4166209102;
        test_addr[7] = 579;
        test_data[7] = 33'd5053671187;
        test_addr[8] = 39;
        test_data[8] = 33'd7928211212;
        test_addr[9] = 345;
        test_data[9] = 33'd2552656500;
        test_addr[10] = 758;
        test_data[10] = 33'd6252825330;
        test_addr[11] = 966;
        test_data[11] = 33'd4123438644;
        test_addr[12] = 994;
        test_data[12] = 33'd2394012061;
        test_addr[13] = 688;
        test_data[13] = 33'd3601440211;
        test_addr[14] = 248;
        test_data[14] = 33'd8455424989;
        test_addr[15] = 466;
        test_data[15] = 33'd3439948819;
        test_addr[16] = 167;
        test_data[16] = 33'd5821482216;
        test_addr[17] = 991;
        test_data[17] = 33'd1186657120;
        test_addr[18] = 371;
        test_data[18] = 33'd2128993578;
        test_addr[19] = 492;
        test_data[19] = 33'd3279720460;
        test_addr[20] = 693;
        test_data[20] = 33'd107943679;
        test_addr[21] = 391;
        test_data[21] = 33'd3059314876;
        test_addr[22] = 3;
        test_data[22] = 33'd2710397198;
        test_addr[23] = 940;
        test_data[23] = 33'd4310782003;
        test_addr[24] = 811;
        test_data[24] = 33'd4521213246;
        test_addr[25] = 180;
        test_data[25] = 33'd1768002488;
        test_addr[26] = 531;
        test_data[26] = 33'd1030173785;
        test_addr[27] = 903;
        test_data[27] = 33'd3268229861;
        test_addr[28] = 714;
        test_data[28] = 33'd4030058467;
        test_addr[29] = 647;
        test_data[29] = 33'd1466466644;
        test_addr[30] = 373;
        test_data[30] = 33'd843400262;
        test_addr[31] = 45;
        test_data[31] = 33'd720913470;
        test_addr[32] = 49;
        test_data[32] = 33'd2053400777;
        test_addr[33] = 375;
        test_data[33] = 33'd116681397;
        test_addr[34] = 32;
        test_data[34] = 33'd7205260702;
        test_addr[35] = 43;
        test_data[35] = 33'd3562471067;
        test_addr[36] = 432;
        test_data[36] = 33'd3643494175;
        test_addr[37] = 358;
        test_data[37] = 33'd6715625422;
        test_addr[38] = 411;
        test_data[38] = 33'd6719221478;
        test_addr[39] = 330;
        test_data[39] = 33'd2270922047;
        test_addr[40] = 319;
        test_data[40] = 33'd7058727247;
        test_addr[41] = 654;
        test_data[41] = 33'd5279750896;
        test_addr[42] = 263;
        test_data[42] = 33'd1115477981;
        test_addr[43] = 136;
        test_data[43] = 33'd933962107;
        test_addr[44] = 684;
        test_data[44] = 33'd4096736423;
        test_addr[45] = 444;
        test_data[45] = 33'd2818036757;
        test_addr[46] = 930;
        test_data[46] = 33'd528430591;
        test_addr[47] = 503;
        test_data[47] = 33'd3936231662;
        test_addr[48] = 961;
        test_data[48] = 33'd5044236111;
        test_addr[49] = 620;
        test_data[49] = 33'd990877164;
        test_addr[50] = 202;
        test_data[50] = 33'd3541495957;
        test_addr[51] = 941;
        test_data[51] = 33'd4153701105;
        test_addr[52] = 31;
        test_data[52] = 33'd2160288399;
        test_addr[53] = 91;
        test_data[53] = 33'd5256460836;
        test_addr[54] = 49;
        test_data[54] = 33'd5736873201;
        test_addr[55] = 484;
        test_data[55] = 33'd3316009856;
        test_addr[56] = 520;
        test_data[56] = 33'd7609894800;
        test_addr[57] = 53;
        test_data[57] = 33'd1440417870;
        test_addr[58] = 879;
        test_data[58] = 33'd978943048;
        test_addr[59] = 281;
        test_data[59] = 33'd8015527480;
        test_addr[60] = 322;
        test_data[60] = 33'd4483009913;
        test_addr[61] = 250;
        test_data[61] = 33'd6472088590;
        test_addr[62] = 755;
        test_data[62] = 33'd1863651176;
        test_addr[63] = 837;
        test_data[63] = 33'd1693487156;
        test_addr[64] = 1003;
        test_data[64] = 33'd8296514786;
        test_addr[65] = 403;
        test_data[65] = 33'd1005991444;
        test_addr[66] = 516;
        test_data[66] = 33'd3801022005;
        test_addr[67] = 597;
        test_data[67] = 33'd2521741564;
        test_addr[68] = 430;
        test_data[68] = 33'd863164190;
        test_addr[69] = 177;
        test_data[69] = 33'd2905827243;
        test_addr[70] = 828;
        test_data[70] = 33'd5402488564;
        test_addr[71] = 613;
        test_data[71] = 33'd1975594517;
        test_addr[72] = 264;
        test_data[72] = 33'd835312204;
        test_addr[73] = 782;
        test_data[73] = 33'd7277731573;
        test_addr[74] = 272;
        test_data[74] = 33'd3167753977;
        test_addr[75] = 970;
        test_data[75] = 33'd3921400631;
        test_addr[76] = 34;
        test_data[76] = 33'd5269658087;
        test_addr[77] = 318;
        test_data[77] = 33'd3083830815;
        test_addr[78] = 803;
        test_data[78] = 33'd3117956401;
        test_addr[79] = 263;
        test_data[79] = 33'd7251859173;
        test_addr[80] = 862;
        test_data[80] = 33'd1375551832;
        test_addr[81] = 637;
        test_data[81] = 33'd2030896509;
        test_addr[82] = 893;
        test_data[82] = 33'd3704026762;
        test_addr[83] = 821;
        test_data[83] = 33'd5234583411;
        test_addr[84] = 920;
        test_data[84] = 33'd1092104427;
        test_addr[85] = 457;
        test_data[85] = 33'd4191839408;
        test_addr[86] = 681;
        test_data[86] = 33'd2735001250;
        test_addr[87] = 206;
        test_data[87] = 33'd7735899550;
        test_addr[88] = 678;
        test_data[88] = 33'd3688685586;
        test_addr[89] = 967;
        test_data[89] = 33'd5992595523;
        test_addr[90] = 370;
        test_data[90] = 33'd4079085858;
        test_addr[91] = 471;
        test_data[91] = 33'd3963935252;
        test_addr[92] = 163;
        test_data[92] = 33'd4051124924;
        test_addr[93] = 486;
        test_data[93] = 33'd4912343941;
        test_addr[94] = 941;
        test_data[94] = 33'd6734675128;
        test_addr[95] = 460;
        test_data[95] = 33'd544566434;
        test_addr[96] = 77;
        test_data[96] = 33'd57221148;
        test_addr[97] = 502;
        test_data[97] = 33'd1213399919;
        test_addr[98] = 220;
        test_data[98] = 33'd1246824563;
        test_addr[99] = 814;
        test_data[99] = 33'd3975966587;
        test_addr[100] = 641;
        test_data[100] = 33'd2076475850;
        test_addr[101] = 46;
        test_data[101] = 33'd2323962822;
        test_addr[102] = 1004;
        test_data[102] = 33'd2043377402;
        test_addr[103] = 533;
        test_data[103] = 33'd5738589063;
        test_addr[104] = 985;
        test_data[104] = 33'd212834635;
        test_addr[105] = 511;
        test_data[105] = 33'd6760035229;
        test_addr[106] = 903;
        test_data[106] = 33'd3268229861;
        test_addr[107] = 615;
        test_data[107] = 33'd3415332789;
        test_addr[108] = 821;
        test_data[108] = 33'd939616115;
        test_addr[109] = 362;
        test_data[109] = 33'd1169309859;
        test_addr[110] = 112;
        test_data[110] = 33'd1757482678;
        test_addr[111] = 113;
        test_data[111] = 33'd419860717;
        test_addr[112] = 22;
        test_data[112] = 33'd2308919392;
        test_addr[113] = 418;
        test_data[113] = 33'd6109325758;
        test_addr[114] = 809;
        test_data[114] = 33'd5494841377;
        test_addr[115] = 346;
        test_data[115] = 33'd4650886467;
        test_addr[116] = 468;
        test_data[116] = 33'd5352947673;
        test_addr[117] = 371;
        test_data[117] = 33'd2128993578;
        test_addr[118] = 64;
        test_data[118] = 33'd1958157960;
        test_addr[119] = 116;
        test_data[119] = 33'd5624203880;
        test_addr[120] = 226;
        test_data[120] = 33'd6427376176;
        test_addr[121] = 25;
        test_data[121] = 33'd6908583646;
        test_addr[122] = 291;
        test_data[122] = 33'd5327708779;
        test_addr[123] = 348;
        test_data[123] = 33'd5762265706;
        test_addr[124] = 327;
        test_data[124] = 33'd614436650;
        test_addr[125] = 466;
        test_data[125] = 33'd3439948819;
        test_addr[126] = 508;
        test_data[126] = 33'd2458412144;
        test_addr[127] = 313;
        test_data[127] = 33'd6515368291;
        test_addr[128] = 639;
        test_data[128] = 33'd3943965978;
        test_addr[129] = 825;
        test_data[129] = 33'd4252998212;
        test_addr[130] = 122;
        test_data[130] = 33'd2514466426;
        test_addr[131] = 500;
        test_data[131] = 33'd8488783149;
        test_addr[132] = 810;
        test_data[132] = 33'd6822723645;
        test_addr[133] = 393;
        test_data[133] = 33'd7322657814;
        test_addr[134] = 655;
        test_data[134] = 33'd300940477;
        test_addr[135] = 23;
        test_data[135] = 33'd2328303965;
        test_addr[136] = 353;
        test_data[136] = 33'd1320710077;
        test_addr[137] = 590;
        test_data[137] = 33'd7816182204;
        test_addr[138] = 66;
        test_data[138] = 33'd1363225947;
        test_addr[139] = 388;
        test_data[139] = 33'd6233848761;
        test_addr[140] = 152;
        test_data[140] = 33'd2706977723;
        test_addr[141] = 444;
        test_data[141] = 33'd2818036757;
        test_addr[142] = 575;
        test_data[142] = 33'd5347607747;
        test_addr[143] = 48;
        test_data[143] = 33'd3954156962;
        test_addr[144] = 948;
        test_data[144] = 33'd2974746974;
        test_addr[145] = 846;
        test_data[145] = 33'd2824502397;
        test_addr[146] = 584;
        test_data[146] = 33'd4559720679;
        test_addr[147] = 52;
        test_data[147] = 33'd3694524907;
        test_addr[148] = 330;
        test_data[148] = 33'd4344530041;
        test_addr[149] = 469;
        test_data[149] = 33'd7963874587;
        test_addr[150] = 899;
        test_data[150] = 33'd5182284847;
        test_addr[151] = 963;
        test_data[151] = 33'd11250872;
        test_addr[152] = 27;
        test_data[152] = 33'd7413626883;
        test_addr[153] = 818;
        test_data[153] = 33'd3235329560;
        test_addr[154] = 168;
        test_data[154] = 33'd8406332547;
        test_addr[155] = 18;
        test_data[155] = 33'd6012427090;
        test_addr[156] = 149;
        test_data[156] = 33'd5624323579;
        test_addr[157] = 921;
        test_data[157] = 33'd2725134890;
        test_addr[158] = 164;
        test_data[158] = 33'd4743396589;
        test_addr[159] = 706;
        test_data[159] = 33'd6415832938;
        test_addr[160] = 317;
        test_data[160] = 33'd7678783066;
        test_addr[161] = 96;
        test_data[161] = 33'd767733627;
        test_addr[162] = 527;
        test_data[162] = 33'd7168663174;
        test_addr[163] = 876;
        test_data[163] = 33'd5662598529;
        test_addr[164] = 97;
        test_data[164] = 33'd62382029;
        test_addr[165] = 851;
        test_data[165] = 33'd1149027704;
        test_addr[166] = 818;
        test_data[166] = 33'd3235329560;
        test_addr[167] = 993;
        test_data[167] = 33'd2081880215;
        test_addr[168] = 576;
        test_data[168] = 33'd4655545476;
        test_addr[169] = 790;
        test_data[169] = 33'd6187296546;
        test_addr[170] = 647;
        test_data[170] = 33'd1466466644;
        test_addr[171] = 641;
        test_data[171] = 33'd2076475850;
        test_addr[172] = 60;
        test_data[172] = 33'd3343706505;
        test_addr[173] = 767;
        test_data[173] = 33'd1189601977;
        test_addr[174] = 679;
        test_data[174] = 33'd2092664236;
        test_addr[175] = 599;
        test_data[175] = 33'd5837394476;
        test_addr[176] = 770;
        test_data[176] = 33'd2171678767;
        test_addr[177] = 581;
        test_data[177] = 33'd1862601448;
        test_addr[178] = 307;
        test_data[178] = 33'd7213693020;
        test_addr[179] = 2;
        test_data[179] = 33'd5154788794;
        test_addr[180] = 506;
        test_data[180] = 33'd659028168;
        test_addr[181] = 296;
        test_data[181] = 33'd5375330532;
        test_addr[182] = 795;
        test_data[182] = 33'd88944858;
        test_addr[183] = 364;
        test_data[183] = 33'd3098727765;
        test_addr[184] = 921;
        test_data[184] = 33'd2725134890;
        test_addr[185] = 42;
        test_data[185] = 33'd4096363574;
        test_addr[186] = 931;
        test_data[186] = 33'd6047340251;
        test_addr[187] = 554;
        test_data[187] = 33'd7817774837;
        test_addr[188] = 21;
        test_data[188] = 33'd789026206;
        test_addr[189] = 854;
        test_data[189] = 33'd8520663752;
        test_addr[190] = 432;
        test_data[190] = 33'd6044307260;
        test_addr[191] = 869;
        test_data[191] = 33'd6106283639;
        test_addr[192] = 262;
        test_data[192] = 33'd7193042145;
        test_addr[193] = 645;
        test_data[193] = 33'd5773575089;
        test_addr[194] = 784;
        test_data[194] = 33'd1428448895;
        test_addr[195] = 496;
        test_data[195] = 33'd8114442729;
        test_addr[196] = 455;
        test_data[196] = 33'd442340444;
        test_addr[197] = 497;
        test_data[197] = 33'd7137838642;
        test_addr[198] = 603;
        test_data[198] = 33'd631643568;
        test_addr[199] = 548;
        test_data[199] = 33'd1224644377;
        test_addr[200] = 827;
        test_data[200] = 33'd6020136494;
        test_addr[201] = 535;
        test_data[201] = 33'd3322326490;
        test_addr[202] = 842;
        test_data[202] = 33'd4586437725;
        test_addr[203] = 506;
        test_data[203] = 33'd659028168;
        test_addr[204] = 208;
        test_data[204] = 33'd881023582;
        test_addr[205] = 500;
        test_data[205] = 33'd4193815853;
        test_addr[206] = 627;
        test_data[206] = 33'd2656035837;
        test_addr[207] = 543;
        test_data[207] = 33'd1828813246;
        test_addr[208] = 423;
        test_data[208] = 33'd6723030281;
        test_addr[209] = 971;
        test_data[209] = 33'd7164180324;
        test_addr[210] = 266;
        test_data[210] = 33'd6773779274;
        test_addr[211] = 703;
        test_data[211] = 33'd3644357459;
        test_addr[212] = 590;
        test_data[212] = 33'd3521214908;
        test_addr[213] = 902;
        test_data[213] = 33'd6779920629;
        test_addr[214] = 446;
        test_data[214] = 33'd1055605986;
        test_addr[215] = 1014;
        test_data[215] = 33'd2402115690;
        test_addr[216] = 889;
        test_data[216] = 33'd3384816046;
        test_addr[217] = 924;
        test_data[217] = 33'd7510846277;
        test_addr[218] = 835;
        test_data[218] = 33'd5346349787;
        test_addr[219] = 166;
        test_data[219] = 33'd6772149917;
        test_addr[220] = 933;
        test_data[220] = 33'd1333871334;
        test_addr[221] = 271;
        test_data[221] = 33'd3753349860;
        test_addr[222] = 389;
        test_data[222] = 33'd7047610350;
        test_addr[223] = 151;
        test_data[223] = 33'd4042063966;
        test_addr[224] = 964;
        test_data[224] = 33'd3846880485;
        test_addr[225] = 725;
        test_data[225] = 33'd7775578593;
        test_addr[226] = 790;
        test_data[226] = 33'd6304902261;
        test_addr[227] = 535;
        test_data[227] = 33'd3322326490;
        test_addr[228] = 123;
        test_data[228] = 33'd3166000446;
        test_addr[229] = 556;
        test_data[229] = 33'd1863958673;
        test_addr[230] = 404;
        test_data[230] = 33'd586528649;
        test_addr[231] = 786;
        test_data[231] = 33'd6645986952;
        test_addr[232] = 93;
        test_data[232] = 33'd7307126697;
        test_addr[233] = 881;
        test_data[233] = 33'd4954896721;
        test_addr[234] = 328;
        test_data[234] = 33'd1334801209;
        test_addr[235] = 713;
        test_data[235] = 33'd358436771;
        test_addr[236] = 742;
        test_data[236] = 33'd4523225485;
        test_addr[237] = 406;
        test_data[237] = 33'd3304677203;
        test_addr[238] = 685;
        test_data[238] = 33'd8500488361;
        test_addr[239] = 69;
        test_data[239] = 33'd445386276;
        test_addr[240] = 448;
        test_data[240] = 33'd6461119132;
        test_addr[241] = 217;
        test_data[241] = 33'd2521597648;
        test_addr[242] = 241;
        test_data[242] = 33'd1993840260;
        test_addr[243] = 514;
        test_data[243] = 33'd1369178089;
        test_addr[244] = 785;
        test_data[244] = 33'd1809300641;
        test_addr[245] = 847;
        test_data[245] = 33'd1925753163;
        test_addr[246] = 459;
        test_data[246] = 33'd8142377452;
        test_addr[247] = 600;
        test_data[247] = 33'd2274691543;
        test_addr[248] = 470;
        test_data[248] = 33'd4198953116;
        test_addr[249] = 590;
        test_data[249] = 33'd3521214908;
        test_addr[250] = 659;
        test_data[250] = 33'd3342857150;
        test_addr[251] = 535;
        test_data[251] = 33'd5222259283;
        test_addr[252] = 962;
        test_data[252] = 33'd1878395484;
        test_addr[253] = 983;
        test_data[253] = 33'd3867328918;
        test_addr[254] = 784;
        test_data[254] = 33'd1428448895;
        test_addr[255] = 59;
        test_data[255] = 33'd1947913714;
        test_addr[256] = 908;
        test_data[256] = 33'd192450639;
        test_addr[257] = 17;
        test_data[257] = 33'd4862448559;
        test_addr[258] = 79;
        test_data[258] = 33'd4243798425;
        test_addr[259] = 892;
        test_data[259] = 33'd2706547949;
        test_addr[260] = 825;
        test_data[260] = 33'd4252998212;
        test_addr[261] = 972;
        test_data[261] = 33'd2852470675;
        test_addr[262] = 419;
        test_data[262] = 33'd4943542373;
        test_addr[263] = 355;
        test_data[263] = 33'd6363863832;
        test_addr[264] = 960;
        test_data[264] = 33'd2916006627;
        test_addr[265] = 329;
        test_data[265] = 33'd7145520034;
        test_addr[266] = 1;
        test_data[266] = 33'd855531051;
        test_addr[267] = 301;
        test_data[267] = 33'd3675695667;
        test_addr[268] = 679;
        test_data[268] = 33'd2092664236;
        test_addr[269] = 123;
        test_data[269] = 33'd3166000446;
        test_addr[270] = 451;
        test_data[270] = 33'd6471461251;
        test_addr[271] = 299;
        test_data[271] = 33'd3042141155;
        test_addr[272] = 635;
        test_data[272] = 33'd7041856570;
        test_addr[273] = 96;
        test_data[273] = 33'd767733627;
        test_addr[274] = 568;
        test_data[274] = 33'd3549289617;
        test_addr[275] = 217;
        test_data[275] = 33'd2521597648;
        test_addr[276] = 214;
        test_data[276] = 33'd6182835276;
        test_addr[277] = 520;
        test_data[277] = 33'd3314927504;
        test_addr[278] = 659;
        test_data[278] = 33'd3342857150;
        test_addr[279] = 49;
        test_data[279] = 33'd5412381996;
        test_addr[280] = 721;
        test_data[280] = 33'd3714234635;
        test_addr[281] = 958;
        test_data[281] = 33'd1861866575;
        test_addr[282] = 655;
        test_data[282] = 33'd7389683545;
        test_addr[283] = 617;
        test_data[283] = 33'd306081816;
        test_addr[284] = 597;
        test_data[284] = 33'd2521741564;
        test_addr[285] = 848;
        test_data[285] = 33'd74868948;
        test_addr[286] = 742;
        test_data[286] = 33'd228258189;
        test_addr[287] = 773;
        test_data[287] = 33'd531933772;
        test_addr[288] = 847;
        test_data[288] = 33'd1925753163;
        test_addr[289] = 156;
        test_data[289] = 33'd7772647361;
        test_addr[290] = 468;
        test_data[290] = 33'd1057980377;
        test_addr[291] = 183;
        test_data[291] = 33'd4082433942;
        test_addr[292] = 490;
        test_data[292] = 33'd309980754;
        test_addr[293] = 564;
        test_data[293] = 33'd1053780301;
        test_addr[294] = 886;
        test_data[294] = 33'd479387173;
        test_addr[295] = 871;
        test_data[295] = 33'd1185961275;
        test_addr[296] = 217;
        test_data[296] = 33'd2521597648;
        test_addr[297] = 511;
        test_data[297] = 33'd2465067933;
        test_addr[298] = 870;
        test_data[298] = 33'd939174474;
        test_addr[299] = 914;
        test_data[299] = 33'd336515192;
        test_addr[300] = 898;
        test_data[300] = 33'd3668671927;
        test_addr[301] = 300;
        test_data[301] = 33'd2360300364;
        test_addr[302] = 570;
        test_data[302] = 33'd1605140899;
        test_addr[303] = 287;
        test_data[303] = 33'd4136431290;
        test_addr[304] = 408;
        test_data[304] = 33'd303432423;
        test_addr[305] = 211;
        test_data[305] = 33'd3319553303;
        test_addr[306] = 1008;
        test_data[306] = 33'd3635208870;
        test_addr[307] = 88;
        test_data[307] = 33'd6341648861;
        test_addr[308] = 967;
        test_data[308] = 33'd1697628227;
        test_addr[309] = 762;
        test_data[309] = 33'd2385791137;
        test_addr[310] = 652;
        test_data[310] = 33'd3031069961;
        test_addr[311] = 797;
        test_data[311] = 33'd3094034019;
        test_addr[312] = 88;
        test_data[312] = 33'd2046681565;
        test_addr[313] = 333;
        test_data[313] = 33'd3264659335;
        test_addr[314] = 300;
        test_data[314] = 33'd2360300364;
        test_addr[315] = 257;
        test_data[315] = 33'd2532794738;
        test_addr[316] = 277;
        test_data[316] = 33'd2128154341;
        test_addr[317] = 619;
        test_data[317] = 33'd3534431847;
        test_addr[318] = 731;
        test_data[318] = 33'd4083566603;
        test_addr[319] = 339;
        test_data[319] = 33'd3510710878;
        test_addr[320] = 263;
        test_data[320] = 33'd2956891877;
        test_addr[321] = 422;
        test_data[321] = 33'd533866239;
        test_addr[322] = 632;
        test_data[322] = 33'd1155677548;
        test_addr[323] = 27;
        test_data[323] = 33'd8526659708;
        test_addr[324] = 512;
        test_data[324] = 33'd3640518258;
        test_addr[325] = 340;
        test_data[325] = 33'd1961019814;
        test_addr[326] = 493;
        test_data[326] = 33'd2901124810;
        test_addr[327] = 1013;
        test_data[327] = 33'd3443847325;
        test_addr[328] = 594;
        test_data[328] = 33'd3713092353;
        test_addr[329] = 60;
        test_data[329] = 33'd5731886175;
        test_addr[330] = 552;
        test_data[330] = 33'd1826755672;
        test_addr[331] = 586;
        test_data[331] = 33'd441018196;
        test_addr[332] = 127;
        test_data[332] = 33'd8051741075;
        test_addr[333] = 856;
        test_data[333] = 33'd4086119564;
        test_addr[334] = 381;
        test_data[334] = 33'd3015459872;
        test_addr[335] = 394;
        test_data[335] = 33'd438437706;
        test_addr[336] = 28;
        test_data[336] = 33'd8174639114;
        test_addr[337] = 185;
        test_data[337] = 33'd4056616662;
        test_addr[338] = 688;
        test_data[338] = 33'd3601440211;
        test_addr[339] = 319;
        test_data[339] = 33'd2763759951;
        test_addr[340] = 285;
        test_data[340] = 33'd705180939;
        test_addr[341] = 180;
        test_data[341] = 33'd5421247094;
        test_addr[342] = 650;
        test_data[342] = 33'd7367325768;
        test_addr[343] = 505;
        test_data[343] = 33'd3673032087;
        test_addr[344] = 823;
        test_data[344] = 33'd700710660;
        test_addr[345] = 777;
        test_data[345] = 33'd850545293;
        test_addr[346] = 717;
        test_data[346] = 33'd3753177976;
        test_addr[347] = 456;
        test_data[347] = 33'd8115338487;
        test_addr[348] = 167;
        test_data[348] = 33'd1526514920;
        test_addr[349] = 224;
        test_data[349] = 33'd643551870;
        test_addr[350] = 733;
        test_data[350] = 33'd1395512612;
        test_addr[351] = 96;
        test_data[351] = 33'd5902467465;
        test_addr[352] = 145;
        test_data[352] = 33'd4495207676;
        test_addr[353] = 920;
        test_data[353] = 33'd1092104427;
        test_addr[354] = 158;
        test_data[354] = 33'd4665608315;
        test_addr[355] = 142;
        test_data[355] = 33'd2263992737;
        test_addr[356] = 980;
        test_data[356] = 33'd5355549282;
        test_addr[357] = 394;
        test_data[357] = 33'd4599416170;
        test_addr[358] = 1023;
        test_data[358] = 33'd107160650;
        test_addr[359] = 441;
        test_data[359] = 33'd948216216;
        test_addr[360] = 698;
        test_data[360] = 33'd3118469034;
        test_addr[361] = 818;
        test_data[361] = 33'd3235329560;
        test_addr[362] = 580;
        test_data[362] = 33'd4090953264;
        test_addr[363] = 504;
        test_data[363] = 33'd3287718623;
        test_addr[364] = 830;
        test_data[364] = 33'd7548746188;
        test_addr[365] = 194;
        test_data[365] = 33'd5369413382;
        test_addr[366] = 288;
        test_data[366] = 33'd262849900;
        test_addr[367] = 351;
        test_data[367] = 33'd7179530918;
        test_addr[368] = 432;
        test_data[368] = 33'd1749339964;
        test_addr[369] = 160;
        test_data[369] = 33'd205033297;
        test_addr[370] = 475;
        test_data[370] = 33'd6853977116;
        test_addr[371] = 1007;
        test_data[371] = 33'd240134872;
        test_addr[372] = 5;
        test_data[372] = 33'd4633374244;
        test_addr[373] = 64;
        test_data[373] = 33'd7307534300;
        test_addr[374] = 439;
        test_data[374] = 33'd3398516884;
        test_addr[375] = 228;
        test_data[375] = 33'd1885599207;
        test_addr[376] = 595;
        test_data[376] = 33'd7500167913;
        test_addr[377] = 787;
        test_data[377] = 33'd2332338642;
        test_addr[378] = 976;
        test_data[378] = 33'd1630561231;
        test_addr[379] = 631;
        test_data[379] = 33'd1893022681;
        test_addr[380] = 830;
        test_data[380] = 33'd3253778892;
        test_addr[381] = 945;
        test_data[381] = 33'd8119400019;
        test_addr[382] = 934;
        test_data[382] = 33'd3429994139;
        test_addr[383] = 741;
        test_data[383] = 33'd1930615449;
        test_addr[384] = 695;
        test_data[384] = 33'd650862610;
        test_addr[385] = 611;
        test_data[385] = 33'd1073177235;
        test_addr[386] = 224;
        test_data[386] = 33'd643551870;
        test_addr[387] = 894;
        test_data[387] = 33'd6587922198;
        test_addr[388] = 930;
        test_data[388] = 33'd6179805919;
        test_addr[389] = 163;
        test_data[389] = 33'd4051124924;
        test_addr[390] = 341;
        test_data[390] = 33'd720341552;
        test_addr[391] = 971;
        test_data[391] = 33'd2869213028;
        test_addr[392] = 30;
        test_data[392] = 33'd561337608;
        test_addr[393] = 811;
        test_data[393] = 33'd226245950;
        test_addr[394] = 93;
        test_data[394] = 33'd3012159401;
        test_addr[395] = 392;
        test_data[395] = 33'd1235012268;
        test_addr[396] = 547;
        test_data[396] = 33'd2078655512;
        test_addr[397] = 221;
        test_data[397] = 33'd2967623187;
        test_addr[398] = 775;
        test_data[398] = 33'd1482893985;
        test_addr[399] = 695;
        test_data[399] = 33'd6289375849;
        test_addr[400] = 7;
        test_data[400] = 33'd2410401329;
        test_addr[401] = 695;
        test_data[401] = 33'd1994408553;
        test_addr[402] = 633;
        test_data[402] = 33'd1648345772;
        test_addr[403] = 244;
        test_data[403] = 33'd2164984734;
        test_addr[404] = 338;
        test_data[404] = 33'd7933654305;
        test_addr[405] = 614;
        test_data[405] = 33'd292281791;
        test_addr[406] = 889;
        test_data[406] = 33'd3384816046;
        test_addr[407] = 397;
        test_data[407] = 33'd7203500539;
        test_addr[408] = 839;
        test_data[408] = 33'd5996659204;
        test_addr[409] = 781;
        test_data[409] = 33'd1625107923;
        test_addr[410] = 922;
        test_data[410] = 33'd3546517031;
        test_addr[411] = 381;
        test_data[411] = 33'd3015459872;
        test_addr[412] = 900;
        test_data[412] = 33'd2793424475;
        test_addr[413] = 326;
        test_data[413] = 33'd6500692716;
        test_addr[414] = 320;
        test_data[414] = 33'd5508035710;
        test_addr[415] = 84;
        test_data[415] = 33'd2985065750;
        test_addr[416] = 860;
        test_data[416] = 33'd5022870474;
        test_addr[417] = 262;
        test_data[417] = 33'd4944359094;
        test_addr[418] = 535;
        test_data[418] = 33'd5998654090;
        test_addr[419] = 687;
        test_data[419] = 33'd6059952363;
        test_addr[420] = 217;
        test_data[420] = 33'd2521597648;
        test_addr[421] = 362;
        test_data[421] = 33'd1169309859;
        test_addr[422] = 492;
        test_data[422] = 33'd8560252878;
        test_addr[423] = 220;
        test_data[423] = 33'd8128390679;
        test_addr[424] = 948;
        test_data[424] = 33'd2974746974;
        test_addr[425] = 941;
        test_data[425] = 33'd8083294857;
        test_addr[426] = 201;
        test_data[426] = 33'd2352154551;
        test_addr[427] = 37;
        test_data[427] = 33'd8408198294;
        test_addr[428] = 172;
        test_data[428] = 33'd1681519392;
        test_addr[429] = 127;
        test_data[429] = 33'd7025459588;
        test_addr[430] = 528;
        test_data[430] = 33'd779927443;
        test_addr[431] = 846;
        test_data[431] = 33'd5870567667;
        test_addr[432] = 542;
        test_data[432] = 33'd5566831229;
        test_addr[433] = 197;
        test_data[433] = 33'd1022834255;
        test_addr[434] = 312;
        test_data[434] = 33'd7888612497;
        test_addr[435] = 60;
        test_data[435] = 33'd1436918879;
        test_addr[436] = 319;
        test_data[436] = 33'd2763759951;
        test_addr[437] = 407;
        test_data[437] = 33'd7832576406;
        test_addr[438] = 132;
        test_data[438] = 33'd438108953;
        test_addr[439] = 94;
        test_data[439] = 33'd4297651294;
        test_addr[440] = 928;
        test_data[440] = 33'd3416090981;
        test_addr[441] = 633;
        test_data[441] = 33'd1648345772;
        test_addr[442] = 182;
        test_data[442] = 33'd3939676421;
        test_addr[443] = 307;
        test_data[443] = 33'd4487592982;
        test_addr[444] = 89;
        test_data[444] = 33'd7907027805;
        test_addr[445] = 307;
        test_data[445] = 33'd192625686;
        test_addr[446] = 904;
        test_data[446] = 33'd4135674155;
        test_addr[447] = 254;
        test_data[447] = 33'd714648240;
        test_addr[448] = 520;
        test_data[448] = 33'd6519200585;
        test_addr[449] = 1011;
        test_data[449] = 33'd5552941075;
        test_addr[450] = 543;
        test_data[450] = 33'd1828813246;
        test_addr[451] = 725;
        test_data[451] = 33'd3480611297;
        test_addr[452] = 172;
        test_data[452] = 33'd1681519392;
        test_addr[453] = 359;
        test_data[453] = 33'd3381025996;
        test_addr[454] = 629;
        test_data[454] = 33'd701803144;
        test_addr[455] = 80;
        test_data[455] = 33'd3551938821;
        test_addr[456] = 156;
        test_data[456] = 33'd3477680065;
        test_addr[457] = 930;
        test_data[457] = 33'd1884838623;
        test_addr[458] = 835;
        test_data[458] = 33'd1051382491;
        test_addr[459] = 178;
        test_data[459] = 33'd3643073190;
        test_addr[460] = 355;
        test_data[460] = 33'd7273705917;
        test_addr[461] = 769;
        test_data[461] = 33'd1388272500;
        test_addr[462] = 189;
        test_data[462] = 33'd2413112707;
        test_addr[463] = 739;
        test_data[463] = 33'd24113143;
        test_addr[464] = 576;
        test_data[464] = 33'd5774271479;
        test_addr[465] = 10;
        test_data[465] = 33'd4272705751;
        test_addr[466] = 792;
        test_data[466] = 33'd758407755;
        test_addr[467] = 793;
        test_data[467] = 33'd7390077616;
        test_addr[468] = 319;
        test_data[468] = 33'd2763759951;
        test_addr[469] = 476;
        test_data[469] = 33'd1210849249;
        test_addr[470] = 491;
        test_data[470] = 33'd1350952293;
        test_addr[471] = 278;
        test_data[471] = 33'd2148021305;
        test_addr[472] = 514;
        test_data[472] = 33'd5643224481;
        test_addr[473] = 412;
        test_data[473] = 33'd38261169;
        test_addr[474] = 595;
        test_data[474] = 33'd7200048739;
        test_addr[475] = 588;
        test_data[475] = 33'd5710177301;
        test_addr[476] = 970;
        test_data[476] = 33'd3921400631;
        test_addr[477] = 188;
        test_data[477] = 33'd3694204641;
        test_addr[478] = 497;
        test_data[478] = 33'd2842871346;
        test_addr[479] = 1018;
        test_data[479] = 33'd1157429103;
        test_addr[480] = 538;
        test_data[480] = 33'd3291868179;
        test_addr[481] = 104;
        test_data[481] = 33'd912554404;
        test_addr[482] = 853;
        test_data[482] = 33'd3949017632;
        test_addr[483] = 76;
        test_data[483] = 33'd1148223066;
        test_addr[484] = 160;
        test_data[484] = 33'd205033297;
        test_addr[485] = 484;
        test_data[485] = 33'd3316009856;
        test_addr[486] = 511;
        test_data[486] = 33'd8371738012;
        test_addr[487] = 271;
        test_data[487] = 33'd3753349860;
        test_addr[488] = 289;
        test_data[488] = 33'd8215964811;
        test_addr[489] = 905;
        test_data[489] = 33'd4369745785;
        test_addr[490] = 934;
        test_data[490] = 33'd4424520922;
        test_addr[491] = 967;
        test_data[491] = 33'd1697628227;
        test_addr[492] = 516;
        test_data[492] = 33'd6059470878;
        test_addr[493] = 394;
        test_data[493] = 33'd304448874;
        test_addr[494] = 212;
        test_data[494] = 33'd51944071;
        test_addr[495] = 92;
        test_data[495] = 33'd11431343;
        test_addr[496] = 403;
        test_data[496] = 33'd7101307036;
        test_addr[497] = 894;
        test_data[497] = 33'd2292954902;
        test_addr[498] = 285;
        test_data[498] = 33'd7530196606;
        test_addr[499] = 121;
        test_data[499] = 33'd8284256091;
        test_addr[500] = 202;
        test_data[500] = 33'd6609565535;
        test_addr[501] = 827;
        test_data[501] = 33'd1725169198;
        test_addr[502] = 363;
        test_data[502] = 33'd3448701357;
        test_addr[503] = 955;
        test_data[503] = 33'd1186627500;
        test_addr[504] = 397;
        test_data[504] = 33'd2908533243;
        test_addr[505] = 685;
        test_data[505] = 33'd6210521411;
        test_addr[506] = 392;
        test_data[506] = 33'd1235012268;
        test_addr[507] = 376;
        test_data[507] = 33'd2751670357;
        test_addr[508] = 1005;
        test_data[508] = 33'd3281370832;
        test_addr[509] = 487;
        test_data[509] = 33'd1196914595;
        test_addr[510] = 585;
        test_data[510] = 33'd7591996435;
        test_addr[511] = 327;
        test_data[511] = 33'd614436650;
        test_addr[512] = 521;
        test_data[512] = 33'd251937582;
        test_addr[513] = 789;
        test_data[513] = 33'd7038325185;
        test_addr[514] = 814;
        test_data[514] = 33'd3975966587;
        test_addr[515] = 137;
        test_data[515] = 33'd6355686352;
        test_addr[516] = 678;
        test_data[516] = 33'd3688685586;
        test_addr[517] = 739;
        test_data[517] = 33'd24113143;
        test_addr[518] = 601;
        test_data[518] = 33'd1792044048;
        test_addr[519] = 376;
        test_data[519] = 33'd2751670357;
        test_addr[520] = 190;
        test_data[520] = 33'd4942286293;
        test_addr[521] = 692;
        test_data[521] = 33'd7776012390;
        test_addr[522] = 792;
        test_data[522] = 33'd758407755;
        test_addr[523] = 35;
        test_data[523] = 33'd3955127962;
        test_addr[524] = 240;
        test_data[524] = 33'd2608724663;
        test_addr[525] = 614;
        test_data[525] = 33'd292281791;
        test_addr[526] = 674;
        test_data[526] = 33'd1833629200;
        test_addr[527] = 937;
        test_data[527] = 33'd7232129049;
        test_addr[528] = 126;
        test_data[528] = 33'd7469058972;
        test_addr[529] = 308;
        test_data[529] = 33'd6599169024;
        test_addr[530] = 653;
        test_data[530] = 33'd7788955784;
        test_addr[531] = 383;
        test_data[531] = 33'd1615749578;
        test_addr[532] = 120;
        test_data[532] = 33'd4431730192;
        test_addr[533] = 997;
        test_data[533] = 33'd7156588838;
        test_addr[534] = 404;
        test_data[534] = 33'd586528649;
        test_addr[535] = 641;
        test_data[535] = 33'd2076475850;
        test_addr[536] = 214;
        test_data[536] = 33'd5572448667;
        test_addr[537] = 768;
        test_data[537] = 33'd7880042411;
        test_addr[538] = 201;
        test_data[538] = 33'd5930463386;
        test_addr[539] = 413;
        test_data[539] = 33'd4791879489;
        test_addr[540] = 50;
        test_data[540] = 33'd6119855017;
        test_addr[541] = 843;
        test_data[541] = 33'd1944986852;
        test_addr[542] = 684;
        test_data[542] = 33'd4096736423;
        test_addr[543] = 772;
        test_data[543] = 33'd925346153;
        test_addr[544] = 814;
        test_data[544] = 33'd6442561713;
        test_addr[545] = 782;
        test_data[545] = 33'd2982764277;
        test_addr[546] = 432;
        test_data[546] = 33'd1749339964;
        test_addr[547] = 106;
        test_data[547] = 33'd7943549416;
        test_addr[548] = 552;
        test_data[548] = 33'd5102278927;
        test_addr[549] = 360;
        test_data[549] = 33'd3720302651;
        test_addr[550] = 464;
        test_data[550] = 33'd1513902136;
        test_addr[551] = 773;
        test_data[551] = 33'd531933772;
        test_addr[552] = 963;
        test_data[552] = 33'd11250872;
        test_addr[553] = 551;
        test_data[553] = 33'd2595070212;
        test_addr[554] = 267;
        test_data[554] = 33'd326083300;
        test_addr[555] = 998;
        test_data[555] = 33'd4165651510;
        test_addr[556] = 478;
        test_data[556] = 33'd2214102913;
        test_addr[557] = 200;
        test_data[557] = 33'd187765645;
        test_addr[558] = 66;
        test_data[558] = 33'd7676754863;
        test_addr[559] = 308;
        test_data[559] = 33'd2304201728;
        test_addr[560] = 520;
        test_data[560] = 33'd2224233289;
        test_addr[561] = 770;
        test_data[561] = 33'd2171678767;
        test_addr[562] = 767;
        test_data[562] = 33'd5952697483;
        test_addr[563] = 689;
        test_data[563] = 33'd753035072;
        test_addr[564] = 533;
        test_data[564] = 33'd6753442654;
        test_addr[565] = 428;
        test_data[565] = 33'd6589693779;
        test_addr[566] = 243;
        test_data[566] = 33'd8315463433;
        test_addr[567] = 596;
        test_data[567] = 33'd1619445656;
        test_addr[568] = 27;
        test_data[568] = 33'd4231692412;
        test_addr[569] = 66;
        test_data[569] = 33'd3381787567;
        test_addr[570] = 95;
        test_data[570] = 33'd4867977810;
        test_addr[571] = 212;
        test_data[571] = 33'd51944071;
        test_addr[572] = 747;
        test_data[572] = 33'd8245496276;
        test_addr[573] = 495;
        test_data[573] = 33'd2224122238;
        test_addr[574] = 881;
        test_data[574] = 33'd6465530667;
        test_addr[575] = 98;
        test_data[575] = 33'd611847547;
        test_addr[576] = 311;
        test_data[576] = 33'd1351719823;
        test_addr[577] = 1013;
        test_data[577] = 33'd3443847325;
        test_addr[578] = 830;
        test_data[578] = 33'd7834241058;
        test_addr[579] = 389;
        test_data[579] = 33'd2752643054;
        test_addr[580] = 656;
        test_data[580] = 33'd2417503440;
        test_addr[581] = 117;
        test_data[581] = 33'd2303502259;
        test_addr[582] = 473;
        test_data[582] = 33'd893693086;
        test_addr[583] = 153;
        test_data[583] = 33'd7740500933;
        test_addr[584] = 905;
        test_data[584] = 33'd8257278787;
        test_addr[585] = 868;
        test_data[585] = 33'd2145195459;
        test_addr[586] = 956;
        test_data[586] = 33'd2021668976;
        test_addr[587] = 954;
        test_data[587] = 33'd643086006;
        test_addr[588] = 980;
        test_data[588] = 33'd1060581986;
        test_addr[589] = 979;
        test_data[589] = 33'd1293811238;
        test_addr[590] = 438;
        test_data[590] = 33'd3272117358;
        test_addr[591] = 908;
        test_data[591] = 33'd192450639;
        test_addr[592] = 64;
        test_data[592] = 33'd3012567004;
        test_addr[593] = 96;
        test_data[593] = 33'd5661514508;
        test_addr[594] = 751;
        test_data[594] = 33'd616267458;
        test_addr[595] = 716;
        test_data[595] = 33'd2231466293;
        test_addr[596] = 878;
        test_data[596] = 33'd1635543175;
        test_addr[597] = 34;
        test_data[597] = 33'd4451512216;
        test_addr[598] = 219;
        test_data[598] = 33'd1413986338;
        test_addr[599] = 622;
        test_data[599] = 33'd981558266;
        test_addr[600] = 132;
        test_data[600] = 33'd438108953;
        test_addr[601] = 585;
        test_data[601] = 33'd7674420448;
        test_addr[602] = 16;
        test_data[602] = 33'd5685208084;
        test_addr[603] = 807;
        test_data[603] = 33'd8557086112;
        test_addr[604] = 757;
        test_data[604] = 33'd1051045639;
        test_addr[605] = 200;
        test_data[605] = 33'd8194768581;
        test_addr[606] = 740;
        test_data[606] = 33'd3140061557;
        test_addr[607] = 403;
        test_data[607] = 33'd6386735609;
        test_addr[608] = 478;
        test_data[608] = 33'd5955056596;
        test_addr[609] = 603;
        test_data[609] = 33'd631643568;
        test_addr[610] = 945;
        test_data[610] = 33'd8202573407;
        test_addr[611] = 1022;
        test_data[611] = 33'd5443014601;
        test_addr[612] = 468;
        test_data[612] = 33'd7913111395;
        test_addr[613] = 499;
        test_data[613] = 33'd3027405431;
        test_addr[614] = 342;
        test_data[614] = 33'd5993354239;
        test_addr[615] = 83;
        test_data[615] = 33'd4027428377;
        test_addr[616] = 116;
        test_data[616] = 33'd1329236584;
        test_addr[617] = 387;
        test_data[617] = 33'd2723287972;
        test_addr[618] = 222;
        test_data[618] = 33'd4085577484;
        test_addr[619] = 657;
        test_data[619] = 33'd927834072;
        test_addr[620] = 1002;
        test_data[620] = 33'd5943041706;
        test_addr[621] = 756;
        test_data[621] = 33'd701769280;
        test_addr[622] = 403;
        test_data[622] = 33'd2091768313;
        test_addr[623] = 829;
        test_data[623] = 33'd1714014072;
        test_addr[624] = 437;
        test_data[624] = 33'd2756765652;
        test_addr[625] = 16;
        test_data[625] = 33'd1390240788;
        test_addr[626] = 516;
        test_data[626] = 33'd1764503582;
        test_addr[627] = 483;
        test_data[627] = 33'd5564248083;
        test_addr[628] = 871;
        test_data[628] = 33'd1185961275;
        test_addr[629] = 1007;
        test_data[629] = 33'd5227095931;
        test_addr[630] = 604;
        test_data[630] = 33'd1821330664;
        test_addr[631] = 352;
        test_data[631] = 33'd4406473444;
        test_addr[632] = 695;
        test_data[632] = 33'd1994408553;
        test_addr[633] = 132;
        test_data[633] = 33'd438108953;
        test_addr[634] = 229;
        test_data[634] = 33'd1480893710;
        test_addr[635] = 974;
        test_data[635] = 33'd4232010606;
        test_addr[636] = 579;
        test_data[636] = 33'd758703891;
        test_addr[637] = 761;
        test_data[637] = 33'd5923111042;
        test_addr[638] = 538;
        test_data[638] = 33'd7389140724;
        test_addr[639] = 58;
        test_data[639] = 33'd6838547580;
        test_addr[640] = 567;
        test_data[640] = 33'd1569593133;
        test_addr[641] = 938;
        test_data[641] = 33'd4486581532;
        test_addr[642] = 521;
        test_data[642] = 33'd251937582;
        test_addr[643] = 442;
        test_data[643] = 33'd5298920770;
        test_addr[644] = 327;
        test_data[644] = 33'd614436650;
        test_addr[645] = 337;
        test_data[645] = 33'd264400746;
        test_addr[646] = 961;
        test_data[646] = 33'd4612378576;
        test_addr[647] = 201;
        test_data[647] = 33'd6054053448;
        test_addr[648] = 597;
        test_data[648] = 33'd2521741564;
        test_addr[649] = 853;
        test_data[649] = 33'd8540060928;
        test_addr[650] = 350;
        test_data[650] = 33'd3916124113;
        test_addr[651] = 459;
        test_data[651] = 33'd3847410156;
        test_addr[652] = 253;
        test_data[652] = 33'd3724959485;
        test_addr[653] = 764;
        test_data[653] = 33'd3790187111;
        test_addr[654] = 715;
        test_data[654] = 33'd662596021;
        test_addr[655] = 436;
        test_data[655] = 33'd3704035340;
        test_addr[656] = 269;
        test_data[656] = 33'd478738172;
        test_addr[657] = 275;
        test_data[657] = 33'd2980684711;
        test_addr[658] = 226;
        test_data[658] = 33'd2132408880;
        test_addr[659] = 332;
        test_data[659] = 33'd5922956456;
        test_addr[660] = 395;
        test_data[660] = 33'd1385063468;
        test_addr[661] = 822;
        test_data[661] = 33'd6685328959;
        test_addr[662] = 562;
        test_data[662] = 33'd3051066239;
        test_addr[663] = 436;
        test_data[663] = 33'd7357044274;
        test_addr[664] = 5;
        test_data[664] = 33'd338406948;
        test_addr[665] = 125;
        test_data[665] = 33'd682282384;
        test_addr[666] = 646;
        test_data[666] = 33'd132734761;
        test_addr[667] = 349;
        test_data[667] = 33'd7151256746;
        test_addr[668] = 82;
        test_data[668] = 33'd2006336925;
        test_addr[669] = 856;
        test_data[669] = 33'd7152544046;
        test_addr[670] = 572;
        test_data[670] = 33'd2425967003;
        test_addr[671] = 298;
        test_data[671] = 33'd6890614106;
        test_addr[672] = 567;
        test_data[672] = 33'd1569593133;
        test_addr[673] = 132;
        test_data[673] = 33'd7445586226;
        test_addr[674] = 377;
        test_data[674] = 33'd4390107465;
        test_addr[675] = 91;
        test_data[675] = 33'd961493540;
        test_addr[676] = 521;
        test_data[676] = 33'd251937582;
        test_addr[677] = 938;
        test_data[677] = 33'd5877341376;
        test_addr[678] = 679;
        test_data[678] = 33'd6405671131;
        test_addr[679] = 749;
        test_data[679] = 33'd1442235455;
        test_addr[680] = 491;
        test_data[680] = 33'd1350952293;
        test_addr[681] = 572;
        test_data[681] = 33'd2425967003;
        test_addr[682] = 46;
        test_data[682] = 33'd5982739849;
        test_addr[683] = 127;
        test_data[683] = 33'd7094346671;
        test_addr[684] = 680;
        test_data[684] = 33'd555640076;
        test_addr[685] = 373;
        test_data[685] = 33'd6039386824;
        test_addr[686] = 107;
        test_data[686] = 33'd5642634824;
        test_addr[687] = 735;
        test_data[687] = 33'd7592571513;
        test_addr[688] = 54;
        test_data[688] = 33'd3762075597;
        test_addr[689] = 173;
        test_data[689] = 33'd2097875581;
        test_addr[690] = 568;
        test_data[690] = 33'd3549289617;
        test_addr[691] = 299;
        test_data[691] = 33'd3042141155;
        test_addr[692] = 979;
        test_data[692] = 33'd1293811238;
        test_addr[693] = 384;
        test_data[693] = 33'd2950368077;
        test_addr[694] = 337;
        test_data[694] = 33'd264400746;
        test_addr[695] = 901;
        test_data[695] = 33'd2235022597;
        test_addr[696] = 126;
        test_data[696] = 33'd3174091676;
        test_addr[697] = 853;
        test_data[697] = 33'd6754726285;
        test_addr[698] = 894;
        test_data[698] = 33'd8283689532;
        test_addr[699] = 603;
        test_data[699] = 33'd631643568;
        test_addr[700] = 442;
        test_data[700] = 33'd1003953474;
        test_addr[701] = 473;
        test_data[701] = 33'd7192831158;
        test_addr[702] = 604;
        test_data[702] = 33'd1821330664;
        test_addr[703] = 38;
        test_data[703] = 33'd1762764931;
        test_addr[704] = 569;
        test_data[704] = 33'd2945905132;
        test_addr[705] = 675;
        test_data[705] = 33'd4804891957;
        test_addr[706] = 871;
        test_data[706] = 33'd1185961275;
        test_addr[707] = 694;
        test_data[707] = 33'd7712055950;
        test_addr[708] = 719;
        test_data[708] = 33'd7698592825;
        test_addr[709] = 922;
        test_data[709] = 33'd3546517031;
        test_addr[710] = 711;
        test_data[710] = 33'd2188493423;
        test_addr[711] = 293;
        test_data[711] = 33'd2329958859;
        test_addr[712] = 122;
        test_data[712] = 33'd4506758699;
        test_addr[713] = 352;
        test_data[713] = 33'd5890784011;
        test_addr[714] = 322;
        test_data[714] = 33'd4925475333;
        test_addr[715] = 559;
        test_data[715] = 33'd4164214068;
        test_addr[716] = 8;
        test_data[716] = 33'd5467897346;
        test_addr[717] = 964;
        test_data[717] = 33'd5767736846;
        test_addr[718] = 531;
        test_data[718] = 33'd5445811369;
        test_addr[719] = 363;
        test_data[719] = 33'd3448701357;
        test_addr[720] = 401;
        test_data[720] = 33'd7738116418;
        test_addr[721] = 88;
        test_data[721] = 33'd2046681565;
        test_addr[722] = 452;
        test_data[722] = 33'd5019387649;
        test_addr[723] = 974;
        test_data[723] = 33'd4232010606;
        test_addr[724] = 882;
        test_data[724] = 33'd1957393229;
        test_addr[725] = 776;
        test_data[725] = 33'd1107570546;
        test_addr[726] = 20;
        test_data[726] = 33'd3947163269;
        test_addr[727] = 987;
        test_data[727] = 33'd4200030814;
        test_addr[728] = 108;
        test_data[728] = 33'd849662807;
        test_addr[729] = 1010;
        test_data[729] = 33'd70305260;
        test_addr[730] = 827;
        test_data[730] = 33'd1725169198;
        test_addr[731] = 404;
        test_data[731] = 33'd586528649;
        test_addr[732] = 152;
        test_data[732] = 33'd4331853581;
        test_addr[733] = 765;
        test_data[733] = 33'd5138819557;
        test_addr[734] = 71;
        test_data[734] = 33'd1938766220;
        test_addr[735] = 341;
        test_data[735] = 33'd720341552;
        test_addr[736] = 921;
        test_data[736] = 33'd2725134890;
        test_addr[737] = 937;
        test_data[737] = 33'd4944971406;
        test_addr[738] = 568;
        test_data[738] = 33'd3549289617;
        test_addr[739] = 283;
        test_data[739] = 33'd3321912760;
        test_addr[740] = 555;
        test_data[740] = 33'd5666177096;
        test_addr[741] = 192;
        test_data[741] = 33'd6015713995;
        test_addr[742] = 186;
        test_data[742] = 33'd3350085156;
        test_addr[743] = 898;
        test_data[743] = 33'd3668671927;
        test_addr[744] = 88;
        test_data[744] = 33'd2046681565;
        test_addr[745] = 1006;
        test_data[745] = 33'd5199787519;
        test_addr[746] = 738;
        test_data[746] = 33'd2491419620;
        test_addr[747] = 79;
        test_data[747] = 33'd4243798425;
        test_addr[748] = 956;
        test_data[748] = 33'd2021668976;
        test_addr[749] = 877;
        test_data[749] = 33'd7901567794;
        test_addr[750] = 2;
        test_data[750] = 33'd859821498;
        test_addr[751] = 666;
        test_data[751] = 33'd1448801851;
        test_addr[752] = 528;
        test_data[752] = 33'd5039686889;
        test_addr[753] = 512;
        test_data[753] = 33'd8505406352;
        test_addr[754] = 915;
        test_data[754] = 33'd275549499;
        test_addr[755] = 697;
        test_data[755] = 33'd8190203451;
        test_addr[756] = 128;
        test_data[756] = 33'd2369463817;
        test_addr[757] = 175;
        test_data[757] = 33'd4616823937;
        test_addr[758] = 232;
        test_data[758] = 33'd4946313757;
        test_addr[759] = 697;
        test_data[759] = 33'd3895236155;
        test_addr[760] = 186;
        test_data[760] = 33'd5977092270;
        test_addr[761] = 523;
        test_data[761] = 33'd662160688;
        test_addr[762] = 584;
        test_data[762] = 33'd264753383;
        test_addr[763] = 446;
        test_data[763] = 33'd1055605986;
        test_addr[764] = 734;
        test_data[764] = 33'd2662220977;
        test_addr[765] = 81;
        test_data[765] = 33'd4489411413;
        test_addr[766] = 526;
        test_data[766] = 33'd512884825;
        test_addr[767] = 619;
        test_data[767] = 33'd3534431847;
        test_addr[768] = 452;
        test_data[768] = 33'd724420353;
        test_addr[769] = 383;
        test_data[769] = 33'd1615749578;
        test_addr[770] = 425;
        test_data[770] = 33'd3413574269;
        test_addr[771] = 996;
        test_data[771] = 33'd3896560801;
        test_addr[772] = 319;
        test_data[772] = 33'd7649728855;
        test_addr[773] = 498;
        test_data[773] = 33'd8005525695;
        test_addr[774] = 151;
        test_data[774] = 33'd4042063966;
        test_addr[775] = 719;
        test_data[775] = 33'd3403625529;
        test_addr[776] = 638;
        test_data[776] = 33'd2536119541;
        test_addr[777] = 530;
        test_data[777] = 33'd3894234752;
        test_addr[778] = 295;
        test_data[778] = 33'd6404470200;
        test_addr[779] = 815;
        test_data[779] = 33'd2868329003;
        test_addr[780] = 64;
        test_data[780] = 33'd5552690849;
        test_addr[781] = 639;
        test_data[781] = 33'd4624581191;
        test_addr[782] = 379;
        test_data[782] = 33'd3734682012;
        test_addr[783] = 106;
        test_data[783] = 33'd4466131988;
        test_addr[784] = 408;
        test_data[784] = 33'd303432423;
        test_addr[785] = 912;
        test_data[785] = 33'd1730083639;
        test_addr[786] = 382;
        test_data[786] = 33'd5001805997;
        test_addr[787] = 731;
        test_data[787] = 33'd5209201607;
        test_addr[788] = 319;
        test_data[788] = 33'd3354761559;
        test_addr[789] = 204;
        test_data[789] = 33'd6811179468;
        test_addr[790] = 603;
        test_data[790] = 33'd6401899771;
        test_addr[791] = 810;
        test_data[791] = 33'd2527756349;
        test_addr[792] = 399;
        test_data[792] = 33'd2238490792;
        test_addr[793] = 380;
        test_data[793] = 33'd4448809795;
        test_addr[794] = 672;
        test_data[794] = 33'd1691338492;
        test_addr[795] = 747;
        test_data[795] = 33'd5196642502;
        test_addr[796] = 954;
        test_data[796] = 33'd643086006;
        test_addr[797] = 191;
        test_data[797] = 33'd3616306016;
        test_addr[798] = 210;
        test_data[798] = 33'd5391219881;
        test_addr[799] = 210;
        test_data[799] = 33'd6425680408;
        test_addr[800] = 815;
        test_data[800] = 33'd8086532860;
        test_addr[801] = 441;
        test_data[801] = 33'd948216216;
        test_addr[802] = 385;
        test_data[802] = 33'd6515740565;
        test_addr[803] = 367;
        test_data[803] = 33'd3102588231;
        test_addr[804] = 274;
        test_data[804] = 33'd3059293611;
        test_addr[805] = 42;
        test_data[805] = 33'd5408577529;
        test_addr[806] = 948;
        test_data[806] = 33'd6361901312;
        test_addr[807] = 1014;
        test_data[807] = 33'd4874928556;
        test_addr[808] = 968;
        test_data[808] = 33'd4989310979;
        test_addr[809] = 418;
        test_data[809] = 33'd1814358462;
        test_addr[810] = 469;
        test_data[810] = 33'd3668907291;
        test_addr[811] = 969;
        test_data[811] = 33'd5888660648;
        test_addr[812] = 712;
        test_data[812] = 33'd3498676098;
        test_addr[813] = 814;
        test_data[813] = 33'd2147594417;
        test_addr[814] = 53;
        test_data[814] = 33'd1440417870;
        test_addr[815] = 101;
        test_data[815] = 33'd334015143;
        test_addr[816] = 194;
        test_data[816] = 33'd1074446086;
        test_addr[817] = 996;
        test_data[817] = 33'd3896560801;
        test_addr[818] = 419;
        test_data[818] = 33'd648575077;
        test_addr[819] = 880;
        test_data[819] = 33'd1460846078;
        test_addr[820] = 798;
        test_data[820] = 33'd8505895484;
        test_addr[821] = 873;
        test_data[821] = 33'd1792266633;
        test_addr[822] = 12;
        test_data[822] = 33'd1981417174;
        test_addr[823] = 384;
        test_data[823] = 33'd6661877969;
        test_addr[824] = 982;
        test_data[824] = 33'd441351460;
        test_addr[825] = 896;
        test_data[825] = 33'd3066857618;
        test_addr[826] = 337;
        test_data[826] = 33'd264400746;
        test_addr[827] = 672;
        test_data[827] = 33'd7753662258;
        test_addr[828] = 683;
        test_data[828] = 33'd3125603621;
        test_addr[829] = 844;
        test_data[829] = 33'd8017462522;
        test_addr[830] = 234;
        test_data[830] = 33'd6798822231;
        test_addr[831] = 622;
        test_data[831] = 33'd981558266;
        test_addr[832] = 618;
        test_data[832] = 33'd2836784331;
        test_addr[833] = 39;
        test_data[833] = 33'd6775480640;
        test_addr[834] = 129;
        test_data[834] = 33'd4027118416;
        test_addr[835] = 216;
        test_data[835] = 33'd3992465811;
        test_addr[836] = 448;
        test_data[836] = 33'd2166151836;
        test_addr[837] = 769;
        test_data[837] = 33'd1388272500;
        test_addr[838] = 745;
        test_data[838] = 33'd2968700236;
        test_addr[839] = 436;
        test_data[839] = 33'd3062076978;
        test_addr[840] = 866;
        test_data[840] = 33'd2280351118;
        test_addr[841] = 578;
        test_data[841] = 33'd5644558338;
        test_addr[842] = 848;
        test_data[842] = 33'd74868948;
        test_addr[843] = 114;
        test_data[843] = 33'd4093300057;
        test_addr[844] = 8;
        test_data[844] = 33'd7409538399;
        test_addr[845] = 53;
        test_data[845] = 33'd8116097155;
        test_addr[846] = 202;
        test_data[846] = 33'd2314598239;
        test_addr[847] = 85;
        test_data[847] = 33'd4465127046;
        test_addr[848] = 517;
        test_data[848] = 33'd4736119378;
        test_addr[849] = 859;
        test_data[849] = 33'd6340410669;
        test_addr[850] = 711;
        test_data[850] = 33'd2188493423;
        test_addr[851] = 73;
        test_data[851] = 33'd261290754;
        test_addr[852] = 1007;
        test_data[852] = 33'd932128635;
        test_addr[853] = 487;
        test_data[853] = 33'd1196914595;
        test_addr[854] = 358;
        test_data[854] = 33'd2420658126;
        test_addr[855] = 533;
        test_data[855] = 33'd6457644551;
        test_addr[856] = 528;
        test_data[856] = 33'd744719593;
        test_addr[857] = 525;
        test_data[857] = 33'd2405063111;
        test_addr[858] = 1007;
        test_data[858] = 33'd932128635;
        test_addr[859] = 843;
        test_data[859] = 33'd4644863909;
        test_addr[860] = 968;
        test_data[860] = 33'd694343683;
        test_addr[861] = 807;
        test_data[861] = 33'd5022426292;
        test_addr[862] = 162;
        test_data[862] = 33'd3110936348;
        test_addr[863] = 161;
        test_data[863] = 33'd5891609294;
        test_addr[864] = 233;
        test_data[864] = 33'd5626152594;
        test_addr[865] = 532;
        test_data[865] = 33'd6794502780;
        test_addr[866] = 621;
        test_data[866] = 33'd7962191918;
        test_addr[867] = 774;
        test_data[867] = 33'd2834186409;
        test_addr[868] = 626;
        test_data[868] = 33'd4427002839;
        test_addr[869] = 646;
        test_data[869] = 33'd132734761;
        test_addr[870] = 358;
        test_data[870] = 33'd2420658126;
        test_addr[871] = 852;
        test_data[871] = 33'd7347549817;
        test_addr[872] = 15;
        test_data[872] = 33'd4529014525;
        test_addr[873] = 873;
        test_data[873] = 33'd1792266633;
        test_addr[874] = 155;
        test_data[874] = 33'd6328501034;
        test_addr[875] = 545;
        test_data[875] = 33'd2528965743;
        test_addr[876] = 231;
        test_data[876] = 33'd660798456;
        test_addr[877] = 203;
        test_data[877] = 33'd1701074922;
        test_addr[878] = 129;
        test_data[878] = 33'd4027118416;
        test_addr[879] = 469;
        test_data[879] = 33'd5289122197;
        test_addr[880] = 519;
        test_data[880] = 33'd4972990633;
        test_addr[881] = 183;
        test_data[881] = 33'd7084223523;
        test_addr[882] = 867;
        test_data[882] = 33'd3206650022;
        test_addr[883] = 939;
        test_data[883] = 33'd3724952086;
        test_addr[884] = 641;
        test_data[884] = 33'd2076475850;
        test_addr[885] = 836;
        test_data[885] = 33'd2452486217;
        test_addr[886] = 45;
        test_data[886] = 33'd5422295311;
        test_addr[887] = 115;
        test_data[887] = 33'd2847575930;
        test_addr[888] = 798;
        test_data[888] = 33'd4210928188;
        test_addr[889] = 949;
        test_data[889] = 33'd4871640285;
        test_addr[890] = 620;
        test_data[890] = 33'd990877164;
        test_addr[891] = 410;
        test_data[891] = 33'd3327850702;
        test_addr[892] = 88;
        test_data[892] = 33'd4438320877;
        test_addr[893] = 525;
        test_data[893] = 33'd7943790721;
        test_addr[894] = 278;
        test_data[894] = 33'd2148021305;
        test_addr[895] = 742;
        test_data[895] = 33'd228258189;
        test_addr[896] = 25;
        test_data[896] = 33'd2613616350;
        test_addr[897] = 826;
        test_data[897] = 33'd7176080038;
        test_addr[898] = 663;
        test_data[898] = 33'd367404024;
        test_addr[899] = 306;
        test_data[899] = 33'd7578475424;
        test_addr[900] = 373;
        test_data[900] = 33'd4302873669;
        test_addr[901] = 432;
        test_data[901] = 33'd5258315185;
        test_addr[902] = 547;
        test_data[902] = 33'd7827222906;
        test_addr[903] = 314;
        test_data[903] = 33'd4198757162;
        test_addr[904] = 972;
        test_data[904] = 33'd2852470675;
        test_addr[905] = 639;
        test_data[905] = 33'd329613895;
        test_addr[906] = 912;
        test_data[906] = 33'd1730083639;
        test_addr[907] = 494;
        test_data[907] = 33'd1860698751;
        test_addr[908] = 287;
        test_data[908] = 33'd4607239598;
        test_addr[909] = 450;
        test_data[909] = 33'd2465959336;
        test_addr[910] = 831;
        test_data[910] = 33'd3525708661;
        test_addr[911] = 997;
        test_data[911] = 33'd8354361230;
        test_addr[912] = 253;
        test_data[912] = 33'd3724959485;
        test_addr[913] = 853;
        test_data[913] = 33'd2459758989;
        test_addr[914] = 94;
        test_data[914] = 33'd2683998;
        test_addr[915] = 833;
        test_data[915] = 33'd2181837440;
        test_addr[916] = 563;
        test_data[916] = 33'd3249157073;
        test_addr[917] = 261;
        test_data[917] = 33'd3806634879;
        test_addr[918] = 28;
        test_data[918] = 33'd5106181386;
        test_addr[919] = 679;
        test_data[919] = 33'd2110703835;
        test_addr[920] = 337;
        test_data[920] = 33'd7850451384;
        test_addr[921] = 208;
        test_data[921] = 33'd881023582;
        test_addr[922] = 902;
        test_data[922] = 33'd4538595075;
        test_addr[923] = 584;
        test_data[923] = 33'd264753383;
        test_addr[924] = 27;
        test_data[924] = 33'd4231692412;
        test_addr[925] = 860;
        test_data[925] = 33'd5144002351;
        test_addr[926] = 621;
        test_data[926] = 33'd3667224622;
        test_addr[927] = 615;
        test_data[927] = 33'd5397688255;
        test_addr[928] = 847;
        test_data[928] = 33'd1925753163;
        test_addr[929] = 788;
        test_data[929] = 33'd3488647823;
        test_addr[930] = 607;
        test_data[930] = 33'd2212965614;
        test_addr[931] = 139;
        test_data[931] = 33'd3271595497;
        test_addr[932] = 223;
        test_data[932] = 33'd3855190456;
        test_addr[933] = 317;
        test_data[933] = 33'd6437004151;
        test_addr[934] = 211;
        test_data[934] = 33'd5189081303;
        test_addr[935] = 277;
        test_data[935] = 33'd7050810898;
        test_addr[936] = 288;
        test_data[936] = 33'd262849900;
        test_addr[937] = 62;
        test_data[937] = 33'd389109591;
        test_addr[938] = 568;
        test_data[938] = 33'd3549289617;
        test_addr[939] = 9;
        test_data[939] = 33'd536276757;
        test_addr[940] = 720;
        test_data[940] = 33'd3049260861;
        test_addr[941] = 818;
        test_data[941] = 33'd3235329560;
        test_addr[942] = 714;
        test_data[942] = 33'd8461492522;
        test_addr[943] = 118;
        test_data[943] = 33'd1346885424;
        test_addr[944] = 119;
        test_data[944] = 33'd3348202238;
        test_addr[945] = 823;
        test_data[945] = 33'd700710660;
        test_addr[946] = 651;
        test_data[946] = 33'd1407051673;
        test_addr[947] = 242;
        test_data[947] = 33'd2171707476;
        test_addr[948] = 394;
        test_data[948] = 33'd304448874;
        test_addr[949] = 27;
        test_data[949] = 33'd4231692412;
        test_addr[950] = 343;
        test_data[950] = 33'd6467097112;
        test_addr[951] = 763;
        test_data[951] = 33'd1119246121;
        test_addr[952] = 194;
        test_data[952] = 33'd1074446086;
        test_addr[953] = 922;
        test_data[953] = 33'd5740464197;
        test_addr[954] = 647;
        test_data[954] = 33'd1466466644;
        test_addr[955] = 118;
        test_data[955] = 33'd4487115284;
        test_addr[956] = 563;
        test_data[956] = 33'd3249157073;
        test_addr[957] = 25;
        test_data[957] = 33'd2613616350;
        test_addr[958] = 207;
        test_data[958] = 33'd5304781843;
        test_addr[959] = 196;
        test_data[959] = 33'd1007003283;
        test_addr[960] = 591;
        test_data[960] = 33'd2185077938;
        test_addr[961] = 680;
        test_data[961] = 33'd6213062561;
        test_addr[962] = 541;
        test_data[962] = 33'd2903716974;
        test_addr[963] = 819;
        test_data[963] = 33'd1751705146;
        test_addr[964] = 657;
        test_data[964] = 33'd927834072;
        test_addr[965] = 743;
        test_data[965] = 33'd4863965533;
        test_addr[966] = 642;
        test_data[966] = 33'd2479303443;
        test_addr[967] = 483;
        test_data[967] = 33'd8363031809;
        test_addr[968] = 294;
        test_data[968] = 33'd4596107355;
        test_addr[969] = 932;
        test_data[969] = 33'd1138021835;
        test_addr[970] = 615;
        test_data[970] = 33'd8566765124;
        test_addr[971] = 741;
        test_data[971] = 33'd1930615449;
        test_addr[972] = 123;
        test_data[972] = 33'd3166000446;
        test_addr[973] = 1012;
        test_data[973] = 33'd3611161271;
        test_addr[974] = 241;
        test_data[974] = 33'd1993840260;
        test_addr[975] = 569;
        test_data[975] = 33'd2945905132;
        test_addr[976] = 604;
        test_data[976] = 33'd1821330664;
        test_addr[977] = 362;
        test_data[977] = 33'd1169309859;
        test_addr[978] = 675;
        test_data[978] = 33'd7929619872;
        test_addr[979] = 650;
        test_data[979] = 33'd3072358472;
        test_addr[980] = 1004;
        test_data[980] = 33'd6276150579;
        test_addr[981] = 261;
        test_data[981] = 33'd3806634879;
        test_addr[982] = 622;
        test_data[982] = 33'd981558266;
        test_addr[983] = 384;
        test_data[983] = 33'd2366910673;
        test_addr[984] = 462;
        test_data[984] = 33'd1029956024;
        test_addr[985] = 997;
        test_data[985] = 33'd7415636435;
        test_addr[986] = 702;
        test_data[986] = 33'd2449747273;
        test_addr[987] = 904;
        test_data[987] = 33'd4135674155;
        test_addr[988] = 531;
        test_data[988] = 33'd1150844073;
        test_addr[989] = 603;
        test_data[989] = 33'd2106932475;
        test_addr[990] = 823;
        test_data[990] = 33'd700710660;
        test_addr[991] = 227;
        test_data[991] = 33'd5237903385;
        test_addr[992] = 789;
        test_data[992] = 33'd2743357889;
        test_addr[993] = 515;
        test_data[993] = 33'd7646879399;
        test_addr[994] = 302;
        test_data[994] = 33'd5390557580;
        test_addr[995] = 964;
        test_data[995] = 33'd1472769550;
        test_addr[996] = 419;
        test_data[996] = 33'd648575077;
        test_addr[997] = 447;
        test_data[997] = 33'd8226526340;
        test_addr[998] = 344;
        test_data[998] = 33'd2140186060;
        test_addr[999] = 176;
        test_data[999] = 33'd5094083564;
        test_addr[1000] = 389;
        test_data[1000] = 33'd2752643054;
        test_addr[1001] = 953;
        test_data[1001] = 33'd6791816372;
        test_addr[1002] = 448;
        test_data[1002] = 33'd2166151836;
        test_addr[1003] = 909;
        test_data[1003] = 33'd1277973101;
        test_addr[1004] = 893;
        test_data[1004] = 33'd8262009820;
        test_addr[1005] = 906;
        test_data[1005] = 33'd3294149566;
        test_addr[1006] = 151;
        test_data[1006] = 33'd4042063966;
        test_addr[1007] = 218;
        test_data[1007] = 33'd4290554056;
        test_addr[1008] = 478;
        test_data[1008] = 33'd4454710708;
        test_addr[1009] = 667;
        test_data[1009] = 33'd3439559431;
        test_addr[1010] = 707;
        test_data[1010] = 33'd1855980571;
        test_addr[1011] = 172;
        test_data[1011] = 33'd5369796678;
        test_addr[1012] = 513;
        test_data[1012] = 33'd2469969087;
        test_addr[1013] = 53;
        test_data[1013] = 33'd8354986908;
        test_addr[1014] = 229;
        test_data[1014] = 33'd1480893710;
        test_addr[1015] = 354;
        test_data[1015] = 33'd1554725479;
        test_addr[1016] = 261;
        test_data[1016] = 33'd3806634879;
        test_addr[1017] = 277;
        test_data[1017] = 33'd2755843602;
        test_addr[1018] = 554;
        test_data[1018] = 33'd6476716051;
        test_addr[1019] = 975;
        test_data[1019] = 33'd3780880889;
        test_addr[1020] = 642;
        test_data[1020] = 33'd7066450600;
        test_addr[1021] = 1002;
        test_data[1021] = 33'd1648074410;
        test_addr[1022] = 504;
        test_data[1022] = 33'd4933935127;
        test_addr[1023] = 709;
        test_data[1023] = 33'd2882321478;
        test_addr[1024] = 577;
        test_data[1024] = 33'd2874325634;
        test_addr[1025] = 233;
        test_data[1025] = 33'd1331185298;
        test_addr[1026] = 89;
        test_data[1026] = 33'd5720247587;
        test_addr[1027] = 495;
        test_data[1027] = 33'd2224122238;
        test_addr[1028] = 184;
        test_data[1028] = 33'd3271992916;
        test_addr[1029] = 431;
        test_data[1029] = 33'd5017071401;
        test_addr[1030] = 808;
        test_data[1030] = 33'd5179413392;
        test_addr[1031] = 348;
        test_data[1031] = 33'd1467298410;
        test_addr[1032] = 202;
        test_data[1032] = 33'd2314598239;
        test_addr[1033] = 138;
        test_data[1033] = 33'd44804164;
        test_addr[1034] = 304;
        test_data[1034] = 33'd885943171;
        test_addr[1035] = 418;
        test_data[1035] = 33'd1814358462;
        test_addr[1036] = 198;
        test_data[1036] = 33'd3924284121;
        test_addr[1037] = 73;
        test_data[1037] = 33'd261290754;
        test_addr[1038] = 510;
        test_data[1038] = 33'd195368792;
        test_addr[1039] = 145;
        test_data[1039] = 33'd200240380;
        test_addr[1040] = 433;
        test_data[1040] = 33'd764669096;
        test_addr[1041] = 863;
        test_data[1041] = 33'd1442050635;
        test_addr[1042] = 809;
        test_data[1042] = 33'd4705643234;
        test_addr[1043] = 64;
        test_data[1043] = 33'd1257723553;
        test_addr[1044] = 455;
        test_data[1044] = 33'd442340444;
        test_addr[1045] = 908;
        test_data[1045] = 33'd7559897362;
        test_addr[1046] = 76;
        test_data[1046] = 33'd1148223066;
        test_addr[1047] = 466;
        test_data[1047] = 33'd6160233983;
        test_addr[1048] = 668;
        test_data[1048] = 33'd1703734548;
        test_addr[1049] = 832;
        test_data[1049] = 33'd8287500940;
        test_addr[1050] = 552;
        test_data[1050] = 33'd807311631;
        test_addr[1051] = 755;
        test_data[1051] = 33'd6360830695;
        test_addr[1052] = 342;
        test_data[1052] = 33'd1698386943;
        test_addr[1053] = 188;
        test_data[1053] = 33'd3694204641;
        test_addr[1054] = 101;
        test_data[1054] = 33'd334015143;
        test_addr[1055] = 208;
        test_data[1055] = 33'd881023582;
        test_addr[1056] = 659;
        test_data[1056] = 33'd7994957662;
        test_addr[1057] = 157;
        test_data[1057] = 33'd7099957097;
        test_addr[1058] = 491;
        test_data[1058] = 33'd8211873232;
        test_addr[1059] = 1016;
        test_data[1059] = 33'd1576676339;
        test_addr[1060] = 576;
        test_data[1060] = 33'd4436488661;
        test_addr[1061] = 407;
        test_data[1061] = 33'd3537609110;
        test_addr[1062] = 301;
        test_data[1062] = 33'd3675695667;
        test_addr[1063] = 553;
        test_data[1063] = 33'd255303072;
        test_addr[1064] = 320;
        test_data[1064] = 33'd1213068414;
        test_addr[1065] = 1009;
        test_data[1065] = 33'd1069602971;
        test_addr[1066] = 305;
        test_data[1066] = 33'd5071011968;
        test_addr[1067] = 850;
        test_data[1067] = 33'd2610616633;
        test_addr[1068] = 390;
        test_data[1068] = 33'd7467997922;
        test_addr[1069] = 963;
        test_data[1069] = 33'd5441603909;
        test_addr[1070] = 651;
        test_data[1070] = 33'd8067785328;
        test_addr[1071] = 560;
        test_data[1071] = 33'd8244117192;
        test_addr[1072] = 96;
        test_data[1072] = 33'd1366547212;
        test_addr[1073] = 724;
        test_data[1073] = 33'd8413184662;
        test_addr[1074] = 25;
        test_data[1074] = 33'd2613616350;
        test_addr[1075] = 558;
        test_data[1075] = 33'd1054185022;
        test_addr[1076] = 824;
        test_data[1076] = 33'd403117584;
        test_addr[1077] = 17;
        test_data[1077] = 33'd567481263;
        test_addr[1078] = 781;
        test_data[1078] = 33'd1625107923;
        test_addr[1079] = 431;
        test_data[1079] = 33'd7012539610;
        test_addr[1080] = 522;
        test_data[1080] = 33'd160969124;
        test_addr[1081] = 94;
        test_data[1081] = 33'd4844306357;
        test_addr[1082] = 894;
        test_data[1082] = 33'd3988722236;
        test_addr[1083] = 115;
        test_data[1083] = 33'd5279806920;
        test_addr[1084] = 945;
        test_data[1084] = 33'd5437151552;
        test_addr[1085] = 958;
        test_data[1085] = 33'd1861866575;
        test_addr[1086] = 976;
        test_data[1086] = 33'd1630561231;
        test_addr[1087] = 799;
        test_data[1087] = 33'd6713925014;
        test_addr[1088] = 20;
        test_data[1088] = 33'd3947163269;
        test_addr[1089] = 624;
        test_data[1089] = 33'd7061718527;
        test_addr[1090] = 256;
        test_data[1090] = 33'd3872731299;
        test_addr[1091] = 432;
        test_data[1091] = 33'd7528300187;
        test_addr[1092] = 660;
        test_data[1092] = 33'd8008078974;
        test_addr[1093] = 1008;
        test_data[1093] = 33'd3635208870;
        test_addr[1094] = 600;
        test_data[1094] = 33'd8022040145;
        test_addr[1095] = 348;
        test_data[1095] = 33'd1467298410;
        test_addr[1096] = 815;
        test_data[1096] = 33'd3791565564;
        test_addr[1097] = 559;
        test_data[1097] = 33'd4482784003;
        test_addr[1098] = 618;
        test_data[1098] = 33'd5480508926;
        test_addr[1099] = 818;
        test_data[1099] = 33'd3235329560;
        test_addr[1100] = 2;
        test_data[1100] = 33'd6643007248;
        test_addr[1101] = 117;
        test_data[1101] = 33'd8021055897;
        test_addr[1102] = 864;
        test_data[1102] = 33'd702666674;
        test_addr[1103] = 247;
        test_data[1103] = 33'd4145441796;
        test_addr[1104] = 126;
        test_data[1104] = 33'd3174091676;
        test_addr[1105] = 886;
        test_data[1105] = 33'd479387173;
        test_addr[1106] = 131;
        test_data[1106] = 33'd3754095223;
        test_addr[1107] = 773;
        test_data[1107] = 33'd531933772;
        test_addr[1108] = 940;
        test_data[1108] = 33'd5527281059;
        test_addr[1109] = 779;
        test_data[1109] = 33'd7531687410;
        test_addr[1110] = 285;
        test_data[1110] = 33'd3235229310;
        test_addr[1111] = 730;
        test_data[1111] = 33'd237210761;
        test_addr[1112] = 403;
        test_data[1112] = 33'd2091768313;
        test_addr[1113] = 522;
        test_data[1113] = 33'd160969124;
        test_addr[1114] = 260;
        test_data[1114] = 33'd2709922654;
        test_addr[1115] = 313;
        test_data[1115] = 33'd2220400995;
        test_addr[1116] = 481;
        test_data[1116] = 33'd1841367641;
        test_addr[1117] = 868;
        test_data[1117] = 33'd2145195459;
        test_addr[1118] = 528;
        test_data[1118] = 33'd744719593;
        test_addr[1119] = 255;
        test_data[1119] = 33'd7432413374;
        test_addr[1120] = 542;
        test_data[1120] = 33'd1271863933;
        test_addr[1121] = 924;
        test_data[1121] = 33'd3215878981;
        test_addr[1122] = 838;
        test_data[1122] = 33'd4110932613;
        test_addr[1123] = 931;
        test_data[1123] = 33'd7683101902;
        test_addr[1124] = 805;
        test_data[1124] = 33'd2845628761;
        test_addr[1125] = 535;
        test_data[1125] = 33'd1703686794;
        test_addr[1126] = 895;
        test_data[1126] = 33'd2712734655;
        test_addr[1127] = 941;
        test_data[1127] = 33'd3788327561;
        test_addr[1128] = 506;
        test_data[1128] = 33'd659028168;
        test_addr[1129] = 645;
        test_data[1129] = 33'd1478607793;
        test_addr[1130] = 111;
        test_data[1130] = 33'd3145322533;
        test_addr[1131] = 532;
        test_data[1131] = 33'd2499535484;
        test_addr[1132] = 549;
        test_data[1132] = 33'd3183535881;
        test_addr[1133] = 537;
        test_data[1133] = 33'd4885500023;
        test_addr[1134] = 699;
        test_data[1134] = 33'd5606680111;
        test_addr[1135] = 806;
        test_data[1135] = 33'd6394163647;
        test_addr[1136] = 947;
        test_data[1136] = 33'd7196308690;
        test_addr[1137] = 845;
        test_data[1137] = 33'd8538310623;
        test_addr[1138] = 545;
        test_data[1138] = 33'd8063223297;
        test_addr[1139] = 315;
        test_data[1139] = 33'd2804730422;
        test_addr[1140] = 463;
        test_data[1140] = 33'd358187220;
        test_addr[1141] = 354;
        test_data[1141] = 33'd1554725479;
        test_addr[1142] = 615;
        test_data[1142] = 33'd4271797828;
        test_addr[1143] = 764;
        test_data[1143] = 33'd3790187111;
        test_addr[1144] = 62;
        test_data[1144] = 33'd389109591;
        test_addr[1145] = 99;
        test_data[1145] = 33'd962759878;
        test_addr[1146] = 560;
        test_data[1146] = 33'd3949149896;
        test_addr[1147] = 203;
        test_data[1147] = 33'd1701074922;
        test_addr[1148] = 213;
        test_data[1148] = 33'd121162192;
        test_addr[1149] = 7;
        test_data[1149] = 33'd2410401329;
        test_addr[1150] = 516;
        test_data[1150] = 33'd1764503582;
        test_addr[1151] = 993;
        test_data[1151] = 33'd2081880215;
        test_addr[1152] = 465;
        test_data[1152] = 33'd4289052588;
        test_addr[1153] = 16;
        test_data[1153] = 33'd1390240788;
        test_addr[1154] = 405;
        test_data[1154] = 33'd3625043014;
        test_addr[1155] = 301;
        test_data[1155] = 33'd3675695667;
        test_addr[1156] = 653;
        test_data[1156] = 33'd8283812473;
        test_addr[1157] = 398;
        test_data[1157] = 33'd5908622380;
        test_addr[1158] = 74;
        test_data[1158] = 33'd8586569289;
        test_addr[1159] = 623;
        test_data[1159] = 33'd1100459140;
        test_addr[1160] = 288;
        test_data[1160] = 33'd262849900;
        test_addr[1161] = 1004;
        test_data[1161] = 33'd1981183283;
        test_addr[1162] = 621;
        test_data[1162] = 33'd3667224622;
        test_addr[1163] = 21;
        test_data[1163] = 33'd789026206;
        test_addr[1164] = 732;
        test_data[1164] = 33'd1612454682;
        test_addr[1165] = 679;
        test_data[1165] = 33'd2110703835;
        test_addr[1166] = 342;
        test_data[1166] = 33'd8017999295;
        test_addr[1167] = 311;
        test_data[1167] = 33'd1351719823;
        test_addr[1168] = 401;
        test_data[1168] = 33'd4899312095;
        test_addr[1169] = 78;
        test_data[1169] = 33'd3865815998;
        test_addr[1170] = 275;
        test_data[1170] = 33'd7525195345;
        test_addr[1171] = 675;
        test_data[1171] = 33'd3634652576;
        test_addr[1172] = 247;
        test_data[1172] = 33'd4145441796;
        test_addr[1173] = 469;
        test_data[1173] = 33'd5743880152;
        test_addr[1174] = 74;
        test_data[1174] = 33'd4291601993;
        test_addr[1175] = 920;
        test_data[1175] = 33'd1092104427;
        test_addr[1176] = 0;
        test_data[1176] = 33'd8480756958;
        test_addr[1177] = 297;
        test_data[1177] = 33'd141773217;
        test_addr[1178] = 945;
        test_data[1178] = 33'd1142184256;
        test_addr[1179] = 752;
        test_data[1179] = 33'd2638568597;
        test_addr[1180] = 899;
        test_data[1180] = 33'd6214310969;
        test_addr[1181] = 469;
        test_data[1181] = 33'd1448912856;
        test_addr[1182] = 184;
        test_data[1182] = 33'd7246230474;
        test_addr[1183] = 847;
        test_data[1183] = 33'd1925753163;
        test_addr[1184] = 54;
        test_data[1184] = 33'd3762075597;
        test_addr[1185] = 209;
        test_data[1185] = 33'd7317197360;
        test_addr[1186] = 394;
        test_data[1186] = 33'd6429176777;
        test_addr[1187] = 478;
        test_data[1187] = 33'd5793520455;
        test_addr[1188] = 740;
        test_data[1188] = 33'd3140061557;
        test_addr[1189] = 315;
        test_data[1189] = 33'd6154387214;
        test_addr[1190] = 252;
        test_data[1190] = 33'd4126756018;
        test_addr[1191] = 837;
        test_data[1191] = 33'd1693487156;
        test_addr[1192] = 829;
        test_data[1192] = 33'd4449865849;
        test_addr[1193] = 472;
        test_data[1193] = 33'd5660774765;
        test_addr[1194] = 704;
        test_data[1194] = 33'd2828619334;
        test_addr[1195] = 375;
        test_data[1195] = 33'd116681397;
        test_addr[1196] = 891;
        test_data[1196] = 33'd2459813267;
        test_addr[1197] = 535;
        test_data[1197] = 33'd4848043120;
        test_addr[1198] = 74;
        test_data[1198] = 33'd6251369512;
        test_addr[1199] = 520;
        test_data[1199] = 33'd2224233289;
        test_addr[1200] = 566;
        test_data[1200] = 33'd3343708057;
        test_addr[1201] = 374;
        test_data[1201] = 33'd7098392497;
        test_addr[1202] = 779;
        test_data[1202] = 33'd3236720114;
        test_addr[1203] = 192;
        test_data[1203] = 33'd1720746699;
        test_addr[1204] = 276;
        test_data[1204] = 33'd5344155853;
        test_addr[1205] = 25;
        test_data[1205] = 33'd2613616350;
        test_addr[1206] = 965;
        test_data[1206] = 33'd2839272030;
        test_addr[1207] = 34;
        test_data[1207] = 33'd6865282830;
        test_addr[1208] = 299;
        test_data[1208] = 33'd3042141155;
        test_addr[1209] = 1003;
        test_data[1209] = 33'd4296035433;
        test_addr[1210] = 931;
        test_data[1210] = 33'd3388134606;
        test_addr[1211] = 405;
        test_data[1211] = 33'd7392686714;
        test_addr[1212] = 360;
        test_data[1212] = 33'd5631144455;
        test_addr[1213] = 1;
        test_data[1213] = 33'd855531051;
        test_addr[1214] = 565;
        test_data[1214] = 33'd8536351826;
        test_addr[1215] = 349;
        test_data[1215] = 33'd4689425632;
        test_addr[1216] = 683;
        test_data[1216] = 33'd6422783047;
        test_addr[1217] = 96;
        test_data[1217] = 33'd1366547212;
        test_addr[1218] = 325;
        test_data[1218] = 33'd3825338226;
        test_addr[1219] = 17;
        test_data[1219] = 33'd567481263;
        test_addr[1220] = 678;
        test_data[1220] = 33'd3688685586;
        test_addr[1221] = 375;
        test_data[1221] = 33'd7865837870;
        test_addr[1222] = 358;
        test_data[1222] = 33'd2420658126;
        test_addr[1223] = 384;
        test_data[1223] = 33'd4842239047;
        test_addr[1224] = 943;
        test_data[1224] = 33'd7017125007;
        test_addr[1225] = 439;
        test_data[1225] = 33'd3398516884;
        test_addr[1226] = 1011;
        test_data[1226] = 33'd1257973779;
        test_addr[1227] = 642;
        test_data[1227] = 33'd2771483304;
        test_addr[1228] = 410;
        test_data[1228] = 33'd7965875563;
        test_addr[1229] = 152;
        test_data[1229] = 33'd36886285;
        test_addr[1230] = 118;
        test_data[1230] = 33'd192147988;
        test_addr[1231] = 1019;
        test_data[1231] = 33'd510091675;
        test_addr[1232] = 652;
        test_data[1232] = 33'd7640163443;
        test_addr[1233] = 285;
        test_data[1233] = 33'd6104402409;
        test_addr[1234] = 256;
        test_data[1234] = 33'd8300044535;
        test_addr[1235] = 397;
        test_data[1235] = 33'd2908533243;
        test_addr[1236] = 988;
        test_data[1236] = 33'd2921234412;
        test_addr[1237] = 529;
        test_data[1237] = 33'd3797362521;
        test_addr[1238] = 975;
        test_data[1238] = 33'd8299719000;
        test_addr[1239] = 677;
        test_data[1239] = 33'd73624117;
        test_addr[1240] = 862;
        test_data[1240] = 33'd7061428402;
        test_addr[1241] = 844;
        test_data[1241] = 33'd6558140893;
        test_addr[1242] = 162;
        test_data[1242] = 33'd3110936348;
        test_addr[1243] = 40;
        test_data[1243] = 33'd3594722951;
        test_addr[1244] = 87;
        test_data[1244] = 33'd3337487982;
        test_addr[1245] = 452;
        test_data[1245] = 33'd6170212670;
        test_addr[1246] = 350;
        test_data[1246] = 33'd6828009009;
        test_addr[1247] = 388;
        test_data[1247] = 33'd1938881465;
        test_addr[1248] = 337;
        test_data[1248] = 33'd3555484088;
        test_addr[1249] = 197;
        test_data[1249] = 33'd1022834255;
        test_addr[1250] = 946;
        test_data[1250] = 33'd8295559936;
        test_addr[1251] = 449;
        test_data[1251] = 33'd3226103403;
        test_addr[1252] = 165;
        test_data[1252] = 33'd190214731;
        test_addr[1253] = 822;
        test_data[1253] = 33'd8221779098;
        test_addr[1254] = 579;
        test_data[1254] = 33'd758703891;
        test_addr[1255] = 182;
        test_data[1255] = 33'd8245702942;
        test_addr[1256] = 976;
        test_data[1256] = 33'd7690720752;
        test_addr[1257] = 817;
        test_data[1257] = 33'd3133004597;
        test_addr[1258] = 600;
        test_data[1258] = 33'd3727072849;
        test_addr[1259] = 775;
        test_data[1259] = 33'd5983762015;
        test_addr[1260] = 770;
        test_data[1260] = 33'd5055053439;
        test_addr[1261] = 506;
        test_data[1261] = 33'd659028168;
        test_addr[1262] = 25;
        test_data[1262] = 33'd5992997963;
        test_addr[1263] = 900;
        test_data[1263] = 33'd2793424475;
        test_addr[1264] = 684;
        test_data[1264] = 33'd4595235005;
        test_addr[1265] = 517;
        test_data[1265] = 33'd441152082;
        test_addr[1266] = 409;
        test_data[1266] = 33'd1379904639;
        test_addr[1267] = 113;
        test_data[1267] = 33'd419860717;
        test_addr[1268] = 607;
        test_data[1268] = 33'd2212965614;
        test_addr[1269] = 255;
        test_data[1269] = 33'd3137446078;
        test_addr[1270] = 1011;
        test_data[1270] = 33'd1257973779;
        test_addr[1271] = 622;
        test_data[1271] = 33'd5299880775;
        test_addr[1272] = 741;
        test_data[1272] = 33'd7255908639;
        test_addr[1273] = 604;
        test_data[1273] = 33'd1821330664;
        test_addr[1274] = 1017;
        test_data[1274] = 33'd770943859;
        test_addr[1275] = 979;
        test_data[1275] = 33'd4468325501;
        test_addr[1276] = 285;
        test_data[1276] = 33'd1809435113;
        test_addr[1277] = 919;
        test_data[1277] = 33'd4037234632;
        test_addr[1278] = 755;
        test_data[1278] = 33'd2065863399;
        test_addr[1279] = 927;
        test_data[1279] = 33'd1780961405;
        test_addr[1280] = 784;
        test_data[1280] = 33'd1428448895;
        test_addr[1281] = 623;
        test_data[1281] = 33'd8501936486;
        test_addr[1282] = 1023;
        test_data[1282] = 33'd107160650;
        test_addr[1283] = 227;
        test_data[1283] = 33'd942936089;
        test_addr[1284] = 675;
        test_data[1284] = 33'd3634652576;
        test_addr[1285] = 555;
        test_data[1285] = 33'd1371209800;
        test_addr[1286] = 971;
        test_data[1286] = 33'd8492495560;
        test_addr[1287] = 153;
        test_data[1287] = 33'd5965141264;
        test_addr[1288] = 428;
        test_data[1288] = 33'd4487858250;
        test_addr[1289] = 700;
        test_data[1289] = 33'd2118661662;
        test_addr[1290] = 288;
        test_data[1290] = 33'd262849900;
        test_addr[1291] = 903;
        test_data[1291] = 33'd3268229861;
        test_addr[1292] = 920;
        test_data[1292] = 33'd1092104427;
        test_addr[1293] = 37;
        test_data[1293] = 33'd5444604736;
        test_addr[1294] = 273;
        test_data[1294] = 33'd2277303350;
        test_addr[1295] = 754;
        test_data[1295] = 33'd2262784563;
        test_addr[1296] = 209;
        test_data[1296] = 33'd3022230064;
        test_addr[1297] = 487;
        test_data[1297] = 33'd1196914595;
        test_addr[1298] = 822;
        test_data[1298] = 33'd8241709677;
        test_addr[1299] = 961;
        test_data[1299] = 33'd317411280;
        test_addr[1300] = 821;
        test_data[1300] = 33'd6626136018;
        test_addr[1301] = 934;
        test_data[1301] = 33'd5330963208;
        test_addr[1302] = 64;
        test_data[1302] = 33'd1257723553;
        test_addr[1303] = 52;
        test_data[1303] = 33'd3694524907;
        test_addr[1304] = 204;
        test_data[1304] = 33'd6852824549;
        test_addr[1305] = 800;
        test_data[1305] = 33'd3860457312;
        test_addr[1306] = 540;
        test_data[1306] = 33'd3411388360;
        test_addr[1307] = 365;
        test_data[1307] = 33'd4037880385;
        test_addr[1308] = 638;
        test_data[1308] = 33'd7114422374;
        test_addr[1309] = 933;
        test_data[1309] = 33'd1333871334;
        test_addr[1310] = 494;
        test_data[1310] = 33'd1860698751;
        test_addr[1311] = 402;
        test_data[1311] = 33'd7142055020;
        test_addr[1312] = 296;
        test_data[1312] = 33'd7478479398;
        test_addr[1313] = 675;
        test_data[1313] = 33'd3634652576;
        test_addr[1314] = 240;
        test_data[1314] = 33'd8361634300;
        test_addr[1315] = 440;
        test_data[1315] = 33'd1696256247;
        test_addr[1316] = 623;
        test_data[1316] = 33'd8571914564;
        test_addr[1317] = 584;
        test_data[1317] = 33'd264753383;
        test_addr[1318] = 873;
        test_data[1318] = 33'd8554636400;
        test_addr[1319] = 815;
        test_data[1319] = 33'd7430927491;
        test_addr[1320] = 901;
        test_data[1320] = 33'd7085812887;
        test_addr[1321] = 183;
        test_data[1321] = 33'd6037162756;
        test_addr[1322] = 766;
        test_data[1322] = 33'd5459190827;
        test_addr[1323] = 292;
        test_data[1323] = 33'd5560828135;
        test_addr[1324] = 828;
        test_data[1324] = 33'd1107521268;
        test_addr[1325] = 502;
        test_data[1325] = 33'd1213399919;
        test_addr[1326] = 946;
        test_data[1326] = 33'd6742785244;
        test_addr[1327] = 102;
        test_data[1327] = 33'd1684138397;
        test_addr[1328] = 857;
        test_data[1328] = 33'd1114468449;
        test_addr[1329] = 254;
        test_data[1329] = 33'd7224865684;
        test_addr[1330] = 664;
        test_data[1330] = 33'd836176777;
        test_addr[1331] = 372;
        test_data[1331] = 33'd1694808878;
        test_addr[1332] = 194;
        test_data[1332] = 33'd1074446086;
        test_addr[1333] = 162;
        test_data[1333] = 33'd6019535544;
        test_addr[1334] = 114;
        test_data[1334] = 33'd7917080067;
        test_addr[1335] = 723;
        test_data[1335] = 33'd2519917846;
        test_addr[1336] = 900;
        test_data[1336] = 33'd2793424475;
        test_addr[1337] = 966;
        test_data[1337] = 33'd4123438644;
        test_addr[1338] = 245;
        test_data[1338] = 33'd8309336303;
        test_addr[1339] = 711;
        test_data[1339] = 33'd8147126720;
        test_addr[1340] = 560;
        test_data[1340] = 33'd4812645315;
        test_addr[1341] = 373;
        test_data[1341] = 33'd7906373;
        test_addr[1342] = 887;
        test_data[1342] = 33'd852431783;
        test_addr[1343] = 779;
        test_data[1343] = 33'd3236720114;
        test_addr[1344] = 418;
        test_data[1344] = 33'd6027906966;
        test_addr[1345] = 946;
        test_data[1345] = 33'd2447817948;
        test_addr[1346] = 905;
        test_data[1346] = 33'd3962311491;
        test_addr[1347] = 697;
        test_data[1347] = 33'd3895236155;
        test_addr[1348] = 420;
        test_data[1348] = 33'd3361591300;
        test_addr[1349] = 17;
        test_data[1349] = 33'd567481263;
        test_addr[1350] = 437;
        test_data[1350] = 33'd7876383461;
        test_addr[1351] = 464;
        test_data[1351] = 33'd1513902136;
        test_addr[1352] = 361;
        test_data[1352] = 33'd3093348283;
        test_addr[1353] = 808;
        test_data[1353] = 33'd884446096;
        test_addr[1354] = 948;
        test_data[1354] = 33'd7803137113;
        test_addr[1355] = 989;
        test_data[1355] = 33'd2993705083;
        test_addr[1356] = 583;
        test_data[1356] = 33'd2629654119;
        test_addr[1357] = 1016;
        test_data[1357] = 33'd1576676339;
        test_addr[1358] = 193;
        test_data[1358] = 33'd1827492103;
        test_addr[1359] = 69;
        test_data[1359] = 33'd445386276;
        test_addr[1360] = 640;
        test_data[1360] = 33'd4932681952;
        test_addr[1361] = 963;
        test_data[1361] = 33'd1146636613;
        test_addr[1362] = 325;
        test_data[1362] = 33'd6254311936;
        test_addr[1363] = 783;
        test_data[1363] = 33'd1379073191;
        test_addr[1364] = 834;
        test_data[1364] = 33'd2481571039;
        test_addr[1365] = 846;
        test_data[1365] = 33'd5153144105;
        test_addr[1366] = 829;
        test_data[1366] = 33'd7060067490;
        test_addr[1367] = 247;
        test_data[1367] = 33'd4870845656;
        test_addr[1368] = 64;
        test_data[1368] = 33'd1257723553;
        test_addr[1369] = 149;
        test_data[1369] = 33'd6563500671;
        test_addr[1370] = 186;
        test_data[1370] = 33'd8040264212;
        test_addr[1371] = 799;
        test_data[1371] = 33'd4737056578;
        test_addr[1372] = 662;
        test_data[1372] = 33'd3196149734;
        test_addr[1373] = 974;
        test_data[1373] = 33'd4232010606;
        test_addr[1374] = 794;
        test_data[1374] = 33'd1845668888;
        test_addr[1375] = 187;
        test_data[1375] = 33'd1241473016;
        test_addr[1376] = 343;
        test_data[1376] = 33'd2172129816;
        test_addr[1377] = 148;
        test_data[1377] = 33'd310279149;
        test_addr[1378] = 526;
        test_data[1378] = 33'd512884825;
        test_addr[1379] = 47;
        test_data[1379] = 33'd5184533518;
        test_addr[1380] = 886;
        test_data[1380] = 33'd479387173;
        test_addr[1381] = 487;
        test_data[1381] = 33'd1196914595;
        test_addr[1382] = 733;
        test_data[1382] = 33'd1395512612;
        test_addr[1383] = 907;
        test_data[1383] = 33'd2677761354;
        test_addr[1384] = 144;
        test_data[1384] = 33'd7711605073;
        test_addr[1385] = 932;
        test_data[1385] = 33'd1138021835;
        test_addr[1386] = 611;
        test_data[1386] = 33'd1073177235;
        test_addr[1387] = 5;
        test_data[1387] = 33'd338406948;
        test_addr[1388] = 468;
        test_data[1388] = 33'd3618144099;
        test_addr[1389] = 931;
        test_data[1389] = 33'd3388134606;
        test_addr[1390] = 93;
        test_data[1390] = 33'd3012159401;
        test_addr[1391] = 622;
        test_data[1391] = 33'd1004913479;
        test_addr[1392] = 1016;
        test_data[1392] = 33'd4295859334;
        test_addr[1393] = 601;
        test_data[1393] = 33'd1792044048;
        test_addr[1394] = 999;
        test_data[1394] = 33'd8183838270;
        test_addr[1395] = 928;
        test_data[1395] = 33'd3416090981;
        test_addr[1396] = 768;
        test_data[1396] = 33'd3585075115;
        test_addr[1397] = 440;
        test_data[1397] = 33'd1696256247;
        test_addr[1398] = 325;
        test_data[1398] = 33'd5483358225;
        test_addr[1399] = 325;
        test_data[1399] = 33'd1188390929;
        test_addr[1400] = 520;
        test_data[1400] = 33'd2224233289;
        test_addr[1401] = 666;
        test_data[1401] = 33'd1448801851;
        test_addr[1402] = 290;
        test_data[1402] = 33'd3259086999;
        test_addr[1403] = 281;
        test_data[1403] = 33'd3720560184;
        test_addr[1404] = 660;
        test_data[1404] = 33'd3713111678;
        test_addr[1405] = 545;
        test_data[1405] = 33'd3768256001;
        test_addr[1406] = 544;
        test_data[1406] = 33'd6803464906;
        test_addr[1407] = 586;
        test_data[1407] = 33'd441018196;
        test_addr[1408] = 324;
        test_data[1408] = 33'd5724077240;
        test_addr[1409] = 502;
        test_data[1409] = 33'd1213399919;
        test_addr[1410] = 476;
        test_data[1410] = 33'd1210849249;
        test_addr[1411] = 51;
        test_data[1411] = 33'd869359556;
        test_addr[1412] = 239;
        test_data[1412] = 33'd948945575;
        test_addr[1413] = 300;
        test_data[1413] = 33'd4460658084;
        test_addr[1414] = 784;
        test_data[1414] = 33'd4534473990;
        test_addr[1415] = 186;
        test_data[1415] = 33'd5928575169;
        test_addr[1416] = 908;
        test_data[1416] = 33'd3264930066;
        test_addr[1417] = 574;
        test_data[1417] = 33'd6825830474;
        test_addr[1418] = 62;
        test_data[1418] = 33'd389109591;
        test_addr[1419] = 96;
        test_data[1419] = 33'd1366547212;
        test_addr[1420] = 129;
        test_data[1420] = 33'd4027118416;
        test_addr[1421] = 314;
        test_data[1421] = 33'd4198757162;
        test_addr[1422] = 532;
        test_data[1422] = 33'd2499535484;
        test_addr[1423] = 362;
        test_data[1423] = 33'd1169309859;
        test_addr[1424] = 308;
        test_data[1424] = 33'd2304201728;
        test_addr[1425] = 725;
        test_data[1425] = 33'd3480611297;
        test_addr[1426] = 1003;
        test_data[1426] = 33'd6165523302;
        test_addr[1427] = 47;
        test_data[1427] = 33'd889566222;
        test_addr[1428] = 785;
        test_data[1428] = 33'd5609492714;
        test_addr[1429] = 717;
        test_data[1429] = 33'd7590501081;
        test_addr[1430] = 644;
        test_data[1430] = 33'd2060679594;
        test_addr[1431] = 533;
        test_data[1431] = 33'd2162677255;
        test_addr[1432] = 704;
        test_data[1432] = 33'd2828619334;
        test_addr[1433] = 542;
        test_data[1433] = 33'd5446371111;
        test_addr[1434] = 490;
        test_data[1434] = 33'd5900709785;
        test_addr[1435] = 124;
        test_data[1435] = 33'd8194474756;
        test_addr[1436] = 430;
        test_data[1436] = 33'd863164190;
        test_addr[1437] = 781;
        test_data[1437] = 33'd1625107923;
        test_addr[1438] = 678;
        test_data[1438] = 33'd3688685586;
        test_addr[1439] = 496;
        test_data[1439] = 33'd3819475433;
        test_addr[1440] = 346;
        test_data[1440] = 33'd355919171;
        test_addr[1441] = 300;
        test_data[1441] = 33'd165690788;
        test_addr[1442] = 989;
        test_data[1442] = 33'd2993705083;
        test_addr[1443] = 667;
        test_data[1443] = 33'd3439559431;
        test_addr[1444] = 116;
        test_data[1444] = 33'd8579125501;
        test_addr[1445] = 772;
        test_data[1445] = 33'd6767882233;
        test_addr[1446] = 457;
        test_data[1446] = 33'd4191839408;
        test_addr[1447] = 515;
        test_data[1447] = 33'd3351912103;
        test_addr[1448] = 594;
        test_data[1448] = 33'd3713092353;
        test_addr[1449] = 624;
        test_data[1449] = 33'd2766751231;
        test_addr[1450] = 156;
        test_data[1450] = 33'd3477680065;
        test_addr[1451] = 658;
        test_data[1451] = 33'd2510800920;
        test_addr[1452] = 515;
        test_data[1452] = 33'd4478277081;
        test_addr[1453] = 835;
        test_data[1453] = 33'd5981814068;
        test_addr[1454] = 537;
        test_data[1454] = 33'd5884000487;
        test_addr[1455] = 859;
        test_data[1455] = 33'd5633416843;
        test_addr[1456] = 523;
        test_data[1456] = 33'd5504192813;
        test_addr[1457] = 154;
        test_data[1457] = 33'd818530140;
        test_addr[1458] = 266;
        test_data[1458] = 33'd2478811978;
        test_addr[1459] = 222;
        test_data[1459] = 33'd7008171226;
        test_addr[1460] = 829;
        test_data[1460] = 33'd6749485816;
        test_addr[1461] = 668;
        test_data[1461] = 33'd4825501314;
        test_addr[1462] = 545;
        test_data[1462] = 33'd7730093254;
        test_addr[1463] = 437;
        test_data[1463] = 33'd3581416165;
        test_addr[1464] = 418;
        test_data[1464] = 33'd1732939670;
        test_addr[1465] = 300;
        test_data[1465] = 33'd5990025906;
        test_addr[1466] = 36;
        test_data[1466] = 33'd4439770930;
        test_addr[1467] = 819;
        test_data[1467] = 33'd6155318973;
        test_addr[1468] = 359;
        test_data[1468] = 33'd3381025996;
        test_addr[1469] = 421;
        test_data[1469] = 33'd8118156320;
        test_addr[1470] = 114;
        test_data[1470] = 33'd3622112771;
        test_addr[1471] = 964;
        test_data[1471] = 33'd4528495732;
        test_addr[1472] = 838;
        test_data[1472] = 33'd4110932613;
        test_addr[1473] = 791;
        test_data[1473] = 33'd1872473622;
        test_addr[1474] = 572;
        test_data[1474] = 33'd2425967003;
        test_addr[1475] = 812;
        test_data[1475] = 33'd2158247624;
        test_addr[1476] = 865;
        test_data[1476] = 33'd6545304978;
        test_addr[1477] = 913;
        test_data[1477] = 33'd81643281;
        test_addr[1478] = 463;
        test_data[1478] = 33'd358187220;
        test_addr[1479] = 635;
        test_data[1479] = 33'd2746889274;
        test_addr[1480] = 321;
        test_data[1480] = 33'd3510587126;
        test_addr[1481] = 574;
        test_data[1481] = 33'd7703600176;
        test_addr[1482] = 564;
        test_data[1482] = 33'd1053780301;
        test_addr[1483] = 169;
        test_data[1483] = 33'd137499134;
        test_addr[1484] = 133;
        test_data[1484] = 33'd2160563348;
        test_addr[1485] = 955;
        test_data[1485] = 33'd1186627500;
        test_addr[1486] = 154;
        test_data[1486] = 33'd818530140;
        test_addr[1487] = 231;
        test_data[1487] = 33'd6866487120;
        test_addr[1488] = 875;
        test_data[1488] = 33'd8575169225;
        test_addr[1489] = 751;
        test_data[1489] = 33'd6481746226;
        test_addr[1490] = 868;
        test_data[1490] = 33'd2145195459;
        test_addr[1491] = 72;
        test_data[1491] = 33'd1907660428;
        test_addr[1492] = 460;
        test_data[1492] = 33'd544566434;
        test_addr[1493] = 846;
        test_data[1493] = 33'd4553201179;
        test_addr[1494] = 62;
        test_data[1494] = 33'd389109591;
        test_addr[1495] = 619;
        test_data[1495] = 33'd5336805652;
        test_addr[1496] = 161;
        test_data[1496] = 33'd1596641998;
        test_addr[1497] = 96;
        test_data[1497] = 33'd1366547212;
        test_addr[1498] = 185;
        test_data[1498] = 33'd7973563340;
        test_addr[1499] = 223;
        test_data[1499] = 33'd3855190456;
        test_addr[1500] = 839;
        test_data[1500] = 33'd1701691908;
        test_addr[1501] = 714;
        test_data[1501] = 33'd4166525226;
        test_addr[1502] = 617;
        test_data[1502] = 33'd306081816;
        test_addr[1503] = 336;
        test_data[1503] = 33'd7226645690;
        test_addr[1504] = 46;
        test_data[1504] = 33'd1687772553;
        test_addr[1505] = 522;
        test_data[1505] = 33'd6350067745;
        test_addr[1506] = 857;
        test_data[1506] = 33'd1114468449;
        test_addr[1507] = 156;
        test_data[1507] = 33'd6380219947;
        test_addr[1508] = 762;
        test_data[1508] = 33'd2385791137;
        test_addr[1509] = 882;
        test_data[1509] = 33'd7010193539;
        test_addr[1510] = 727;
        test_data[1510] = 33'd2548078876;
        test_addr[1511] = 103;
        test_data[1511] = 33'd3519285150;
        test_addr[1512] = 434;
        test_data[1512] = 33'd425295928;
        test_addr[1513] = 958;
        test_data[1513] = 33'd8365140169;
        test_addr[1514] = 593;
        test_data[1514] = 33'd4289367533;
        test_addr[1515] = 188;
        test_data[1515] = 33'd6899042248;
        test_addr[1516] = 373;
        test_data[1516] = 33'd7906373;
        test_addr[1517] = 987;
        test_data[1517] = 33'd4200030814;
        test_addr[1518] = 1017;
        test_data[1518] = 33'd770943859;
        test_addr[1519] = 324;
        test_data[1519] = 33'd5574666391;
        test_addr[1520] = 653;
        test_data[1520] = 33'd7969835682;
        test_addr[1521] = 426;
        test_data[1521] = 33'd5863838786;
        test_addr[1522] = 119;
        test_data[1522] = 33'd3348202238;
        test_addr[1523] = 745;
        test_data[1523] = 33'd2968700236;
        test_addr[1524] = 42;
        test_data[1524] = 33'd1113610233;
        test_addr[1525] = 576;
        test_data[1525] = 33'd7816129174;
        test_addr[1526] = 416;
        test_data[1526] = 33'd593392457;
        test_addr[1527] = 835;
        test_data[1527] = 33'd1686846772;
        test_addr[1528] = 438;
        test_data[1528] = 33'd3272117358;
        test_addr[1529] = 48;
        test_data[1529] = 33'd3954156962;
        test_addr[1530] = 713;
        test_data[1530] = 33'd358436771;
        test_addr[1531] = 900;
        test_data[1531] = 33'd2793424475;
        test_addr[1532] = 228;
        test_data[1532] = 33'd1885599207;
        test_addr[1533] = 306;
        test_data[1533] = 33'd3283508128;
        test_addr[1534] = 183;
        test_data[1534] = 33'd1742195460;
        test_addr[1535] = 836;
        test_data[1535] = 33'd2452486217;
        test_addr[1536] = 772;
        test_data[1536] = 33'd2472914937;
        test_addr[1537] = 914;
        test_data[1537] = 33'd336515192;
        test_addr[1538] = 791;
        test_data[1538] = 33'd7567275627;
        test_addr[1539] = 327;
        test_data[1539] = 33'd614436650;
        test_addr[1540] = 466;
        test_data[1540] = 33'd4400496053;
        test_addr[1541] = 979;
        test_data[1541] = 33'd173358205;
        test_addr[1542] = 958;
        test_data[1542] = 33'd4070172873;
        test_addr[1543] = 251;
        test_data[1543] = 33'd7379802526;
        test_addr[1544] = 720;
        test_data[1544] = 33'd3049260861;
        test_addr[1545] = 776;
        test_data[1545] = 33'd1107570546;
        test_addr[1546] = 582;
        test_data[1546] = 33'd3203865679;
        test_addr[1547] = 575;
        test_data[1547] = 33'd8381006396;
        test_addr[1548] = 511;
        test_data[1548] = 33'd4076770716;
        test_addr[1549] = 691;
        test_data[1549] = 33'd3704402127;
        test_addr[1550] = 530;
        test_data[1550] = 33'd6861790606;
        test_addr[1551] = 932;
        test_data[1551] = 33'd6137741236;
        test_addr[1552] = 772;
        test_data[1552] = 33'd7502407474;
        test_addr[1553] = 25;
        test_data[1553] = 33'd1698030667;
        test_addr[1554] = 157;
        test_data[1554] = 33'd2804989801;
        test_addr[1555] = 245;
        test_data[1555] = 33'd5661507185;
        test_addr[1556] = 386;
        test_data[1556] = 33'd1528358932;
        test_addr[1557] = 699;
        test_data[1557] = 33'd7845842621;
        test_addr[1558] = 764;
        test_data[1558] = 33'd3790187111;
        test_addr[1559] = 149;
        test_data[1559] = 33'd4391451060;
        test_addr[1560] = 365;
        test_data[1560] = 33'd7703829080;
        test_addr[1561] = 290;
        test_data[1561] = 33'd3259086999;
        test_addr[1562] = 61;
        test_data[1562] = 33'd3050866392;
        test_addr[1563] = 885;
        test_data[1563] = 33'd8377754463;
        test_addr[1564] = 40;
        test_data[1564] = 33'd3594722951;
        test_addr[1565] = 180;
        test_data[1565] = 33'd1126279798;
        test_addr[1566] = 38;
        test_data[1566] = 33'd1762764931;
        test_addr[1567] = 886;
        test_data[1567] = 33'd479387173;
        test_addr[1568] = 543;
        test_data[1568] = 33'd5887816566;
        test_addr[1569] = 46;
        test_data[1569] = 33'd1687772553;
        test_addr[1570] = 424;
        test_data[1570] = 33'd1637986519;
        test_addr[1571] = 947;
        test_data[1571] = 33'd2901341394;
        test_addr[1572] = 415;
        test_data[1572] = 33'd4390712257;
        test_addr[1573] = 423;
        test_data[1573] = 33'd2428062985;
        test_addr[1574] = 631;
        test_data[1574] = 33'd1893022681;
        test_addr[1575] = 234;
        test_data[1575] = 33'd4576094175;
        test_addr[1576] = 163;
        test_data[1576] = 33'd7962408818;
        test_addr[1577] = 708;
        test_data[1577] = 33'd4183077687;
        test_addr[1578] = 298;
        test_data[1578] = 33'd2595646810;
        test_addr[1579] = 467;
        test_data[1579] = 33'd3833684444;
        test_addr[1580] = 915;
        test_data[1580] = 33'd5288824777;
        test_addr[1581] = 909;
        test_data[1581] = 33'd7359575432;
        test_addr[1582] = 205;
        test_data[1582] = 33'd7478063952;
        test_addr[1583] = 637;
        test_data[1583] = 33'd2030896509;
        test_addr[1584] = 236;
        test_data[1584] = 33'd3976153366;
        test_addr[1585] = 51;
        test_data[1585] = 33'd4860727649;
        test_addr[1586] = 728;
        test_data[1586] = 33'd820874592;
        test_addr[1587] = 286;
        test_data[1587] = 33'd667168271;
        test_addr[1588] = 123;
        test_data[1588] = 33'd4365089074;
        test_addr[1589] = 71;
        test_data[1589] = 33'd1938766220;
        test_addr[1590] = 459;
        test_data[1590] = 33'd5256044891;
        test_addr[1591] = 641;
        test_data[1591] = 33'd2076475850;
        test_addr[1592] = 105;
        test_data[1592] = 33'd1192418195;
        test_addr[1593] = 776;
        test_data[1593] = 33'd6704830763;
        test_addr[1594] = 197;
        test_data[1594] = 33'd1022834255;
        test_addr[1595] = 686;
        test_data[1595] = 33'd4286094390;
        test_addr[1596] = 679;
        test_data[1596] = 33'd2110703835;
        test_addr[1597] = 14;
        test_data[1597] = 33'd7295927927;
        test_addr[1598] = 990;
        test_data[1598] = 33'd616895957;
        test_addr[1599] = 327;
        test_data[1599] = 33'd6603553455;
        test_addr[1600] = 375;
        test_data[1600] = 33'd3570870574;
        test_addr[1601] = 704;
        test_data[1601] = 33'd2828619334;
        test_addr[1602] = 432;
        test_data[1602] = 33'd3233332891;
        test_addr[1603] = 302;
        test_data[1603] = 33'd1095590284;
        test_addr[1604] = 18;
        test_data[1604] = 33'd1717459794;
        test_addr[1605] = 613;
        test_data[1605] = 33'd1975594517;
        test_addr[1606] = 717;
        test_data[1606] = 33'd7019863191;
        test_addr[1607] = 930;
        test_data[1607] = 33'd7133161359;
        test_addr[1608] = 534;
        test_data[1608] = 33'd8287325302;
        test_addr[1609] = 982;
        test_data[1609] = 33'd441351460;
        test_addr[1610] = 166;
        test_data[1610] = 33'd7715315760;
        test_addr[1611] = 135;
        test_data[1611] = 33'd3089281077;
        test_addr[1612] = 441;
        test_data[1612] = 33'd948216216;
        test_addr[1613] = 685;
        test_data[1613] = 33'd7290562329;
        test_addr[1614] = 737;
        test_data[1614] = 33'd1797063890;
        test_addr[1615] = 250;
        test_data[1615] = 33'd6419947008;
        test_addr[1616] = 467;
        test_data[1616] = 33'd3833684444;
        test_addr[1617] = 668;
        test_data[1617] = 33'd530534018;
        test_addr[1618] = 623;
        test_data[1618] = 33'd4276947268;
        test_addr[1619] = 934;
        test_data[1619] = 33'd1035995912;
        test_addr[1620] = 203;
        test_data[1620] = 33'd1701074922;
        test_addr[1621] = 966;
        test_data[1621] = 33'd4123438644;
        test_addr[1622] = 6;
        test_data[1622] = 33'd5723525347;
        test_addr[1623] = 574;
        test_data[1623] = 33'd7683417466;
        test_addr[1624] = 85;
        test_data[1624] = 33'd4369987674;
        test_addr[1625] = 269;
        test_data[1625] = 33'd478738172;
        test_addr[1626] = 653;
        test_data[1626] = 33'd3674868386;
        test_addr[1627] = 217;
        test_data[1627] = 33'd2521597648;
        test_addr[1628] = 1022;
        test_data[1628] = 33'd1148047305;
        test_addr[1629] = 183;
        test_data[1629] = 33'd4299410139;
        test_addr[1630] = 891;
        test_data[1630] = 33'd6153161126;
        test_addr[1631] = 902;
        test_data[1631] = 33'd5537067467;
        test_addr[1632] = 747;
        test_data[1632] = 33'd901675206;
        test_addr[1633] = 932;
        test_data[1633] = 33'd1842773940;
        test_addr[1634] = 715;
        test_data[1634] = 33'd8403692523;
        test_addr[1635] = 449;
        test_data[1635] = 33'd3226103403;
        test_addr[1636] = 645;
        test_data[1636] = 33'd1478607793;
        test_addr[1637] = 723;
        test_data[1637] = 33'd2519917846;
        test_addr[1638] = 769;
        test_data[1638] = 33'd7406167242;
        test_addr[1639] = 512;
        test_data[1639] = 33'd4210439056;
        test_addr[1640] = 938;
        test_data[1640] = 33'd5914085791;
        test_addr[1641] = 167;
        test_data[1641] = 33'd7728870399;
        test_addr[1642] = 837;
        test_data[1642] = 33'd1693487156;
        test_addr[1643] = 847;
        test_data[1643] = 33'd1925753163;
        test_addr[1644] = 618;
        test_data[1644] = 33'd5345096157;
        test_addr[1645] = 284;
        test_data[1645] = 33'd258676554;
        test_addr[1646] = 893;
        test_data[1646] = 33'd3967042524;
        test_addr[1647] = 1000;
        test_data[1647] = 33'd3122678110;
        test_addr[1648] = 552;
        test_data[1648] = 33'd807311631;
        test_addr[1649] = 87;
        test_data[1649] = 33'd7685547776;
        test_addr[1650] = 757;
        test_data[1650] = 33'd1051045639;
        test_addr[1651] = 60;
        test_data[1651] = 33'd1436918879;
        test_addr[1652] = 830;
        test_data[1652] = 33'd3539273762;
        test_addr[1653] = 411;
        test_data[1653] = 33'd2424254182;
        test_addr[1654] = 622;
        test_data[1654] = 33'd1004913479;
        test_addr[1655] = 515;
        test_data[1655] = 33'd183309785;
        test_addr[1656] = 461;
        test_data[1656] = 33'd2300259007;
        test_addr[1657] = 488;
        test_data[1657] = 33'd5488331317;
        test_addr[1658] = 491;
        test_data[1658] = 33'd4812784179;
        test_addr[1659] = 528;
        test_data[1659] = 33'd7199522862;
        test_addr[1660] = 728;
        test_data[1660] = 33'd820874592;
        test_addr[1661] = 532;
        test_data[1661] = 33'd2499535484;
        test_addr[1662] = 808;
        test_data[1662] = 33'd884446096;
        test_addr[1663] = 666;
        test_data[1663] = 33'd1448801851;
        test_addr[1664] = 345;
        test_data[1664] = 33'd5376265032;
        test_addr[1665] = 856;
        test_data[1665] = 33'd2857576750;
        test_addr[1666] = 498;
        test_data[1666] = 33'd3710558399;
        test_addr[1667] = 580;
        test_data[1667] = 33'd4090953264;
        test_addr[1668] = 710;
        test_data[1668] = 33'd7599695076;
        test_addr[1669] = 233;
        test_data[1669] = 33'd1331185298;
        test_addr[1670] = 938;
        test_data[1670] = 33'd4348452935;
        test_addr[1671] = 897;
        test_data[1671] = 33'd1039575909;
        test_addr[1672] = 458;
        test_data[1672] = 33'd6273378637;
        test_addr[1673] = 934;
        test_data[1673] = 33'd1035995912;
        test_addr[1674] = 635;
        test_data[1674] = 33'd7360809762;
        test_addr[1675] = 160;
        test_data[1675] = 33'd205033297;
        test_addr[1676] = 224;
        test_data[1676] = 33'd643551870;
        test_addr[1677] = 779;
        test_data[1677] = 33'd3236720114;
        test_addr[1678] = 224;
        test_data[1678] = 33'd6533024272;
        test_addr[1679] = 541;
        test_data[1679] = 33'd2903716974;
        test_addr[1680] = 114;
        test_data[1680] = 33'd3622112771;
        test_addr[1681] = 968;
        test_data[1681] = 33'd8143337727;
        test_addr[1682] = 76;
        test_data[1682] = 33'd4943756399;
        test_addr[1683] = 27;
        test_data[1683] = 33'd5503978352;
        test_addr[1684] = 29;
        test_data[1684] = 33'd4050089466;
        test_addr[1685] = 352;
        test_data[1685] = 33'd1595816715;
        test_addr[1686] = 56;
        test_data[1686] = 33'd5740675352;
        test_addr[1687] = 456;
        test_data[1687] = 33'd3820371191;
        test_addr[1688] = 747;
        test_data[1688] = 33'd901675206;
        test_addr[1689] = 466;
        test_data[1689] = 33'd105528757;
        test_addr[1690] = 509;
        test_data[1690] = 33'd2005844869;
        test_addr[1691] = 846;
        test_data[1691] = 33'd258233883;
        test_addr[1692] = 843;
        test_data[1692] = 33'd5631367323;
        test_addr[1693] = 91;
        test_data[1693] = 33'd961493540;
        test_addr[1694] = 509;
        test_data[1694] = 33'd2005844869;
        test_addr[1695] = 857;
        test_data[1695] = 33'd1114468449;
        test_addr[1696] = 262;
        test_data[1696] = 33'd649391798;
        test_addr[1697] = 407;
        test_data[1697] = 33'd3537609110;
        test_addr[1698] = 479;
        test_data[1698] = 33'd6615117692;
        test_addr[1699] = 299;
        test_data[1699] = 33'd3042141155;
        test_addr[1700] = 430;
        test_data[1700] = 33'd863164190;
        test_addr[1701] = 453;
        test_data[1701] = 33'd3500901833;
        test_addr[1702] = 258;
        test_data[1702] = 33'd1832274105;
        test_addr[1703] = 445;
        test_data[1703] = 33'd495816375;
        test_addr[1704] = 639;
        test_data[1704] = 33'd329613895;
        test_addr[1705] = 866;
        test_data[1705] = 33'd2280351118;
        test_addr[1706] = 178;
        test_data[1706] = 33'd8002976532;
        test_addr[1707] = 495;
        test_data[1707] = 33'd2224122238;
        test_addr[1708] = 718;
        test_data[1708] = 33'd5446496977;
        test_addr[1709] = 193;
        test_data[1709] = 33'd1827492103;
        test_addr[1710] = 831;
        test_data[1710] = 33'd6681673590;
        test_addr[1711] = 270;
        test_data[1711] = 33'd8312223369;
        test_addr[1712] = 693;
        test_data[1712] = 33'd107943679;
        test_addr[1713] = 730;
        test_data[1713] = 33'd4338827055;
        test_addr[1714] = 100;
        test_data[1714] = 33'd6475816011;
        test_addr[1715] = 101;
        test_data[1715] = 33'd334015143;
        test_addr[1716] = 154;
        test_data[1716] = 33'd818530140;
        test_addr[1717] = 307;
        test_data[1717] = 33'd192625686;
        test_addr[1718] = 20;
        test_data[1718] = 33'd3947163269;
        test_addr[1719] = 617;
        test_data[1719] = 33'd306081816;
        test_addr[1720] = 957;
        test_data[1720] = 33'd1537653831;
        test_addr[1721] = 259;
        test_data[1721] = 33'd1475111032;
        test_addr[1722] = 318;
        test_data[1722] = 33'd6867488296;
        test_addr[1723] = 472;
        test_data[1723] = 33'd1365807469;
        test_addr[1724] = 599;
        test_data[1724] = 33'd1542427180;
        test_addr[1725] = 64;
        test_data[1725] = 33'd1257723553;
        test_addr[1726] = 913;
        test_data[1726] = 33'd81643281;
        test_addr[1727] = 31;
        test_data[1727] = 33'd2160288399;
        test_addr[1728] = 253;
        test_data[1728] = 33'd3724959485;
        test_addr[1729] = 698;
        test_data[1729] = 33'd3118469034;
        test_addr[1730] = 594;
        test_data[1730] = 33'd3713092353;
        test_addr[1731] = 371;
        test_data[1731] = 33'd5063821176;
        test_addr[1732] = 193;
        test_data[1732] = 33'd7890194095;
        test_addr[1733] = 348;
        test_data[1733] = 33'd8216305540;
        test_addr[1734] = 962;
        test_data[1734] = 33'd1878395484;
        test_addr[1735] = 354;
        test_data[1735] = 33'd1554725479;
        test_addr[1736] = 785;
        test_data[1736] = 33'd4823830749;
        test_addr[1737] = 810;
        test_data[1737] = 33'd4315297191;
        test_addr[1738] = 214;
        test_data[1738] = 33'd1277481371;
        test_addr[1739] = 460;
        test_data[1739] = 33'd544566434;
        test_addr[1740] = 670;
        test_data[1740] = 33'd5269375;
        test_addr[1741] = 875;
        test_data[1741] = 33'd6783351898;
        test_addr[1742] = 421;
        test_data[1742] = 33'd6170831325;
        test_addr[1743] = 764;
        test_data[1743] = 33'd3790187111;
        test_addr[1744] = 1001;
        test_data[1744] = 33'd2446236361;
        test_addr[1745] = 773;
        test_data[1745] = 33'd531933772;
        test_addr[1746] = 186;
        test_data[1746] = 33'd8345860302;
        test_addr[1747] = 1004;
        test_data[1747] = 33'd1981183283;
        test_addr[1748] = 478;
        test_data[1748] = 33'd7093890323;
        test_addr[1749] = 552;
        test_data[1749] = 33'd807311631;
        test_addr[1750] = 343;
        test_data[1750] = 33'd2172129816;
        test_addr[1751] = 402;
        test_data[1751] = 33'd2847087724;
        test_addr[1752] = 876;
        test_data[1752] = 33'd5517880342;
        test_addr[1753] = 275;
        test_data[1753] = 33'd8174373852;
        test_addr[1754] = 994;
        test_data[1754] = 33'd2394012061;
        test_addr[1755] = 708;
        test_data[1755] = 33'd4183077687;
        test_addr[1756] = 908;
        test_data[1756] = 33'd3264930066;
        test_addr[1757] = 916;
        test_data[1757] = 33'd379022188;
        test_addr[1758] = 69;
        test_data[1758] = 33'd445386276;
        test_addr[1759] = 354;
        test_data[1759] = 33'd1554725479;
        test_addr[1760] = 533;
        test_data[1760] = 33'd2162677255;
        test_addr[1761] = 228;
        test_data[1761] = 33'd1885599207;
        test_addr[1762] = 220;
        test_data[1762] = 33'd3833423383;
        test_addr[1763] = 996;
        test_data[1763] = 33'd3896560801;
        test_addr[1764] = 852;
        test_data[1764] = 33'd7980282749;
        test_addr[1765] = 859;
        test_data[1765] = 33'd1338449547;
        test_addr[1766] = 645;
        test_data[1766] = 33'd1478607793;
        test_addr[1767] = 4;
        test_data[1767] = 33'd5438707178;
        test_addr[1768] = 19;
        test_data[1768] = 33'd2697384543;
        test_addr[1769] = 530;
        test_data[1769] = 33'd7778419790;
        test_addr[1770] = 866;
        test_data[1770] = 33'd6914695043;
        test_addr[1771] = 656;
        test_data[1771] = 33'd8481173335;
        test_addr[1772] = 467;
        test_data[1772] = 33'd3833684444;
        test_addr[1773] = 757;
        test_data[1773] = 33'd1051045639;
        test_addr[1774] = 655;
        test_data[1774] = 33'd3094716249;
        test_addr[1775] = 342;
        test_data[1775] = 33'd6270473909;
        test_addr[1776] = 74;
        test_data[1776] = 33'd1956402216;
        test_addr[1777] = 267;
        test_data[1777] = 33'd5199745084;
        test_addr[1778] = 720;
        test_data[1778] = 33'd5579279390;
        test_addr[1779] = 735;
        test_data[1779] = 33'd3297604217;
        test_addr[1780] = 379;
        test_data[1780] = 33'd3734682012;
        test_addr[1781] = 813;
        test_data[1781] = 33'd7469747854;
        test_addr[1782] = 237;
        test_data[1782] = 33'd5739678170;
        test_addr[1783] = 786;
        test_data[1783] = 33'd2351019656;
        test_addr[1784] = 659;
        test_data[1784] = 33'd3699990366;
        test_addr[1785] = 995;
        test_data[1785] = 33'd6140114967;
        test_addr[1786] = 314;
        test_data[1786] = 33'd5443243292;
        test_addr[1787] = 289;
        test_data[1787] = 33'd3920997515;
        test_addr[1788] = 238;
        test_data[1788] = 33'd83366238;
        test_addr[1789] = 232;
        test_data[1789] = 33'd5461135377;
        test_addr[1790] = 491;
        test_data[1790] = 33'd517816883;
        test_addr[1791] = 21;
        test_data[1791] = 33'd789026206;
        test_addr[1792] = 884;
        test_data[1792] = 33'd678817658;
        test_addr[1793] = 545;
        test_data[1793] = 33'd6938135033;
        test_addr[1794] = 487;
        test_data[1794] = 33'd1196914595;
        test_addr[1795] = 588;
        test_data[1795] = 33'd1415210005;
        test_addr[1796] = 314;
        test_data[1796] = 33'd1148275996;
        test_addr[1797] = 867;
        test_data[1797] = 33'd6289006749;
        test_addr[1798] = 192;
        test_data[1798] = 33'd5035365690;
        test_addr[1799] = 13;
        test_data[1799] = 33'd7511479614;
        test_addr[1800] = 109;
        test_data[1800] = 33'd2687315092;
        test_addr[1801] = 129;
        test_data[1801] = 33'd7633881987;
        test_addr[1802] = 841;
        test_data[1802] = 33'd7154894208;
        test_addr[1803] = 81;
        test_data[1803] = 33'd4856584088;
        test_addr[1804] = 783;
        test_data[1804] = 33'd1379073191;
        test_addr[1805] = 759;
        test_data[1805] = 33'd2171230616;
        test_addr[1806] = 242;
        test_data[1806] = 33'd2171707476;
        test_addr[1807] = 423;
        test_data[1807] = 33'd2428062985;
        test_addr[1808] = 689;
        test_data[1808] = 33'd753035072;
        test_addr[1809] = 617;
        test_data[1809] = 33'd306081816;
        test_addr[1810] = 105;
        test_data[1810] = 33'd1192418195;
        test_addr[1811] = 207;
        test_data[1811] = 33'd8563566793;
        test_addr[1812] = 462;
        test_data[1812] = 33'd1029956024;
        test_addr[1813] = 127;
        test_data[1813] = 33'd2799379375;
        test_addr[1814] = 379;
        test_data[1814] = 33'd3734682012;
        test_addr[1815] = 794;
        test_data[1815] = 33'd1845668888;
        test_addr[1816] = 448;
        test_data[1816] = 33'd2166151836;
        test_addr[1817] = 900;
        test_data[1817] = 33'd2793424475;
        test_addr[1818] = 431;
        test_data[1818] = 33'd2717572314;
        test_addr[1819] = 813;
        test_data[1819] = 33'd3174780558;
        test_addr[1820] = 970;
        test_data[1820] = 33'd3921400631;
        test_addr[1821] = 49;
        test_data[1821] = 33'd1117414700;
        test_addr[1822] = 381;
        test_data[1822] = 33'd3015459872;
        test_addr[1823] = 642;
        test_data[1823] = 33'd2771483304;
        test_addr[1824] = 82;
        test_data[1824] = 33'd2006336925;
        test_addr[1825] = 752;
        test_data[1825] = 33'd7422541163;
        test_addr[1826] = 609;
        test_data[1826] = 33'd779641857;
        test_addr[1827] = 687;
        test_data[1827] = 33'd6627436173;
        test_addr[1828] = 420;
        test_data[1828] = 33'd3361591300;
        test_addr[1829] = 862;
        test_data[1829] = 33'd5594246134;
        test_addr[1830] = 303;
        test_data[1830] = 33'd3582560146;
        test_addr[1831] = 317;
        test_data[1831] = 33'd2142036855;
        test_addr[1832] = 480;
        test_data[1832] = 33'd2118543923;
        test_addr[1833] = 926;
        test_data[1833] = 33'd2655641510;
        test_addr[1834] = 170;
        test_data[1834] = 33'd1650688480;
        test_addr[1835] = 670;
        test_data[1835] = 33'd5269375;
        test_addr[1836] = 256;
        test_data[1836] = 33'd4005077239;
        test_addr[1837] = 984;
        test_data[1837] = 33'd2904690682;
        test_addr[1838] = 361;
        test_data[1838] = 33'd5585022349;
        test_addr[1839] = 859;
        test_data[1839] = 33'd1338449547;
        test_addr[1840] = 80;
        test_data[1840] = 33'd3551938821;
        test_addr[1841] = 971;
        test_data[1841] = 33'd4197528264;
        test_addr[1842] = 868;
        test_data[1842] = 33'd2145195459;
        test_addr[1843] = 546;
        test_data[1843] = 33'd3391432801;
        test_addr[1844] = 380;
        test_data[1844] = 33'd6555048600;
        test_addr[1845] = 321;
        test_data[1845] = 33'd3510587126;
        test_addr[1846] = 473;
        test_data[1846] = 33'd2897863862;
        test_addr[1847] = 741;
        test_data[1847] = 33'd2960941343;
        test_addr[1848] = 464;
        test_data[1848] = 33'd8054210437;
        test_addr[1849] = 429;
        test_data[1849] = 33'd1861495304;
        test_addr[1850] = 316;
        test_data[1850] = 33'd8326157606;
        test_addr[1851] = 803;
        test_data[1851] = 33'd3117956401;
        test_addr[1852] = 749;
        test_data[1852] = 33'd1442235455;
        test_addr[1853] = 16;
        test_data[1853] = 33'd1390240788;
        test_addr[1854] = 783;
        test_data[1854] = 33'd1379073191;
        test_addr[1855] = 172;
        test_data[1855] = 33'd7823017477;
        test_addr[1856] = 890;
        test_data[1856] = 33'd1732209976;
        test_addr[1857] = 852;
        test_data[1857] = 33'd3685315453;
        test_addr[1858] = 465;
        test_data[1858] = 33'd4289052588;
        test_addr[1859] = 872;
        test_data[1859] = 33'd1431148747;
        test_addr[1860] = 381;
        test_data[1860] = 33'd3015459872;
        test_addr[1861] = 807;
        test_data[1861] = 33'd727458996;
        test_addr[1862] = 137;
        test_data[1862] = 33'd8235606630;
        test_addr[1863] = 82;
        test_data[1863] = 33'd2006336925;
        test_addr[1864] = 837;
        test_data[1864] = 33'd1693487156;
        test_addr[1865] = 340;
        test_data[1865] = 33'd7945645541;
        test_addr[1866] = 166;
        test_data[1866] = 33'd3420348464;
        test_addr[1867] = 440;
        test_data[1867] = 33'd5084171152;
        test_addr[1868] = 197;
        test_data[1868] = 33'd8438761844;
        test_addr[1869] = 591;
        test_data[1869] = 33'd2185077938;
        test_addr[1870] = 937;
        test_data[1870] = 33'd650004110;
        test_addr[1871] = 8;
        test_data[1871] = 33'd3114571103;
        test_addr[1872] = 987;
        test_data[1872] = 33'd8011084240;
        test_addr[1873] = 595;
        test_data[1873] = 33'd2905081443;
        test_addr[1874] = 818;
        test_data[1874] = 33'd6224891476;
        test_addr[1875] = 692;
        test_data[1875] = 33'd3481045094;
        test_addr[1876] = 596;
        test_data[1876] = 33'd1619445656;
        test_addr[1877] = 390;
        test_data[1877] = 33'd7119297222;
        test_addr[1878] = 861;
        test_data[1878] = 33'd3560847281;
        test_addr[1879] = 89;
        test_data[1879] = 33'd1425280291;
        test_addr[1880] = 436;
        test_data[1880] = 33'd3062076978;
        test_addr[1881] = 118;
        test_data[1881] = 33'd192147988;
        test_addr[1882] = 829;
        test_data[1882] = 33'd2454518520;
        test_addr[1883] = 633;
        test_data[1883] = 33'd1648345772;
        test_addr[1884] = 417;
        test_data[1884] = 33'd6900760489;
        test_addr[1885] = 42;
        test_data[1885] = 33'd1113610233;
        test_addr[1886] = 823;
        test_data[1886] = 33'd700710660;
        test_addr[1887] = 810;
        test_data[1887] = 33'd7957854742;
        test_addr[1888] = 385;
        test_data[1888] = 33'd2220773269;
        test_addr[1889] = 636;
        test_data[1889] = 33'd4864859791;
        test_addr[1890] = 550;
        test_data[1890] = 33'd5799212174;
        test_addr[1891] = 216;
        test_data[1891] = 33'd3992465811;
        test_addr[1892] = 970;
        test_data[1892] = 33'd4497261481;
        test_addr[1893] = 803;
        test_data[1893] = 33'd4417544979;
        test_addr[1894] = 351;
        test_data[1894] = 33'd8327940489;
        test_addr[1895] = 25;
        test_data[1895] = 33'd1698030667;
        test_addr[1896] = 148;
        test_data[1896] = 33'd310279149;
        test_addr[1897] = 837;
        test_data[1897] = 33'd1693487156;
        test_addr[1898] = 441;
        test_data[1898] = 33'd948216216;
        test_addr[1899] = 685;
        test_data[1899] = 33'd2995595033;
        test_addr[1900] = 160;
        test_data[1900] = 33'd205033297;
        test_addr[1901] = 412;
        test_data[1901] = 33'd7132834895;
        test_addr[1902] = 675;
        test_data[1902] = 33'd7295736522;
        test_addr[1903] = 29;
        test_data[1903] = 33'd5550253222;
        test_addr[1904] = 415;
        test_data[1904] = 33'd95744961;
        test_addr[1905] = 270;
        test_data[1905] = 33'd6940387313;
        test_addr[1906] = 974;
        test_data[1906] = 33'd4232010606;
        test_addr[1907] = 372;
        test_data[1907] = 33'd1694808878;
        test_addr[1908] = 705;
        test_data[1908] = 33'd3595301892;
        test_addr[1909] = 395;
        test_data[1909] = 33'd1385063468;
        test_addr[1910] = 974;
        test_data[1910] = 33'd7774894007;
        test_addr[1911] = 966;
        test_data[1911] = 33'd4123438644;
        test_addr[1912] = 174;
        test_data[1912] = 33'd7885104970;
        test_addr[1913] = 393;
        test_data[1913] = 33'd4550908162;
        test_addr[1914] = 636;
        test_data[1914] = 33'd6149267026;
        test_addr[1915] = 878;
        test_data[1915] = 33'd1635543175;
        test_addr[1916] = 298;
        test_data[1916] = 33'd2595646810;
        test_addr[1917] = 476;
        test_data[1917] = 33'd1210849249;
        test_addr[1918] = 729;
        test_data[1918] = 33'd1893345796;
        test_addr[1919] = 401;
        test_data[1919] = 33'd6087894323;
        test_addr[1920] = 156;
        test_data[1920] = 33'd6450569423;
        test_addr[1921] = 157;
        test_data[1921] = 33'd8441551675;
        test_addr[1922] = 472;
        test_data[1922] = 33'd1365807469;
        test_addr[1923] = 0;
        test_data[1923] = 33'd7372261257;
        test_addr[1924] = 813;
        test_data[1924] = 33'd3174780558;
        test_addr[1925] = 994;
        test_data[1925] = 33'd4944877549;
        test_addr[1926] = 491;
        test_data[1926] = 33'd517816883;
        test_addr[1927] = 765;
        test_data[1927] = 33'd843852261;
        test_addr[1928] = 705;
        test_data[1928] = 33'd3595301892;
        test_addr[1929] = 509;
        test_data[1929] = 33'd2005844869;
        test_addr[1930] = 789;
        test_data[1930] = 33'd2743357889;
        test_addr[1931] = 971;
        test_data[1931] = 33'd4197528264;
        test_addr[1932] = 638;
        test_data[1932] = 33'd6719158449;
        test_addr[1933] = 860;
        test_data[1933] = 33'd849035055;
        test_addr[1934] = 215;
        test_data[1934] = 33'd815101909;
        test_addr[1935] = 837;
        test_data[1935] = 33'd1693487156;
        test_addr[1936] = 433;
        test_data[1936] = 33'd764669096;
        test_addr[1937] = 741;
        test_data[1937] = 33'd5142487982;
        test_addr[1938] = 690;
        test_data[1938] = 33'd4288616562;
        test_addr[1939] = 813;
        test_data[1939] = 33'd4838466454;
        test_addr[1940] = 709;
        test_data[1940] = 33'd6388945029;
        test_addr[1941] = 546;
        test_data[1941] = 33'd3391432801;
        test_addr[1942] = 7;
        test_data[1942] = 33'd6618079911;
        test_addr[1943] = 860;
        test_data[1943] = 33'd4857733372;
        test_addr[1944] = 13;
        test_data[1944] = 33'd3216512318;
        test_addr[1945] = 872;
        test_data[1945] = 33'd1431148747;
        test_addr[1946] = 322;
        test_data[1946] = 33'd4320974869;
        test_addr[1947] = 401;
        test_data[1947] = 33'd1792927027;
        test_addr[1948] = 715;
        test_data[1948] = 33'd4108725227;
        test_addr[1949] = 803;
        test_data[1949] = 33'd122577683;
        test_addr[1950] = 897;
        test_data[1950] = 33'd1039575909;
        test_addr[1951] = 927;
        test_data[1951] = 33'd1780961405;
        test_addr[1952] = 528;
        test_data[1952] = 33'd2904555566;
        test_addr[1953] = 877;
        test_data[1953] = 33'd3606600498;
        test_addr[1954] = 995;
        test_data[1954] = 33'd7929931471;
        test_addr[1955] = 1012;
        test_data[1955] = 33'd3611161271;
        test_addr[1956] = 949;
        test_data[1956] = 33'd7496737913;
        test_addr[1957] = 737;
        test_data[1957] = 33'd1797063890;
        test_addr[1958] = 756;
        test_data[1958] = 33'd701769280;
        test_addr[1959] = 184;
        test_data[1959] = 33'd2951263178;
        test_addr[1960] = 619;
        test_data[1960] = 33'd1041838356;
        test_addr[1961] = 553;
        test_data[1961] = 33'd255303072;
        test_addr[1962] = 80;
        test_data[1962] = 33'd3551938821;
        test_addr[1963] = 54;
        test_data[1963] = 33'd3762075597;
        test_addr[1964] = 651;
        test_data[1964] = 33'd3772818032;
        test_addr[1965] = 360;
        test_data[1965] = 33'd1336177159;
        test_addr[1966] = 858;
        test_data[1966] = 33'd1864704728;
        test_addr[1967] = 622;
        test_data[1967] = 33'd8292558942;
        test_addr[1968] = 706;
        test_data[1968] = 33'd2120865642;
        test_addr[1969] = 352;
        test_data[1969] = 33'd1595816715;
        test_addr[1970] = 591;
        test_data[1970] = 33'd2185077938;
        test_addr[1971] = 594;
        test_data[1971] = 33'd4511066996;
        test_addr[1972] = 472;
        test_data[1972] = 33'd5089632236;
        test_addr[1973] = 507;
        test_data[1973] = 33'd3886571279;
        test_addr[1974] = 724;
        test_data[1974] = 33'd4118217366;
        test_addr[1975] = 953;
        test_data[1975] = 33'd2496849076;
        test_addr[1976] = 937;
        test_data[1976] = 33'd650004110;
        test_addr[1977] = 773;
        test_data[1977] = 33'd531933772;
        test_addr[1978] = 690;
        test_data[1978] = 33'd4288616562;
        test_addr[1979] = 219;
        test_data[1979] = 33'd6556723714;
        test_addr[1980] = 51;
        test_data[1980] = 33'd565760353;
        test_addr[1981] = 331;
        test_data[1981] = 33'd2402963099;
        test_addr[1982] = 455;
        test_data[1982] = 33'd8455966777;
        test_addr[1983] = 426;
        test_data[1983] = 33'd1568871490;
        test_addr[1984] = 372;
        test_data[1984] = 33'd1694808878;
        test_addr[1985] = 456;
        test_data[1985] = 33'd3820371191;
        test_addr[1986] = 176;
        test_data[1986] = 33'd799116268;
        test_addr[1987] = 513;
        test_data[1987] = 33'd2469969087;
        test_addr[1988] = 1009;
        test_data[1988] = 33'd8234822696;
        test_addr[1989] = 993;
        test_data[1989] = 33'd7460091032;
        test_addr[1990] = 998;
        test_data[1990] = 33'd4165651510;
        test_addr[1991] = 293;
        test_data[1991] = 33'd2329958859;
        test_addr[1992] = 521;
        test_data[1992] = 33'd4848288352;
        test_addr[1993] = 89;
        test_data[1993] = 33'd1425280291;
        test_addr[1994] = 597;
        test_data[1994] = 33'd2521741564;
        test_addr[1995] = 885;
        test_data[1995] = 33'd4082787167;
        test_addr[1996] = 599;
        test_data[1996] = 33'd1542427180;
        test_addr[1997] = 434;
        test_data[1997] = 33'd4473266731;
        test_addr[1998] = 496;
        test_data[1998] = 33'd4557845274;
        test_addr[1999] = 811;
        test_data[1999] = 33'd226245950;
        test_addr[2000] = 255;
        test_data[2000] = 33'd3137446078;
        test_addr[2001] = 865;
        test_data[2001] = 33'd8395913018;
        test_addr[2002] = 414;
        test_data[2002] = 33'd998493570;
        test_addr[2003] = 32;
        test_data[2003] = 33'd4561908415;
        test_addr[2004] = 216;
        test_data[2004] = 33'd6161222379;
        test_addr[2005] = 977;
        test_data[2005] = 33'd4221183128;
        test_addr[2006] = 151;
        test_data[2006] = 33'd4042063966;
        test_addr[2007] = 470;
        test_data[2007] = 33'd4198953116;
        test_addr[2008] = 986;
        test_data[2008] = 33'd942798349;
        test_addr[2009] = 831;
        test_data[2009] = 33'd2386706294;
        test_addr[2010] = 68;
        test_data[2010] = 33'd780007243;
        test_addr[2011] = 195;
        test_data[2011] = 33'd2074235098;
        test_addr[2012] = 588;
        test_data[2012] = 33'd4892175615;
        test_addr[2013] = 666;
        test_data[2013] = 33'd6247440514;
        test_addr[2014] = 465;
        test_data[2014] = 33'd4289052588;
        test_addr[2015] = 260;
        test_data[2015] = 33'd2709922654;
        test_addr[2016] = 782;
        test_data[2016] = 33'd2982764277;
        test_addr[2017] = 257;
        test_data[2017] = 33'd6594620398;
        test_addr[2018] = 908;
        test_data[2018] = 33'd7388570798;
        test_addr[2019] = 536;
        test_data[2019] = 33'd1287154060;
        test_addr[2020] = 492;
        test_data[2020] = 33'd4265285582;
        test_addr[2021] = 861;
        test_data[2021] = 33'd3560847281;
        test_addr[2022] = 895;
        test_data[2022] = 33'd2712734655;
        test_addr[2023] = 587;
        test_data[2023] = 33'd7875651109;
        test_addr[2024] = 569;
        test_data[2024] = 33'd6927986738;
        test_addr[2025] = 446;
        test_data[2025] = 33'd1055605986;
        test_addr[2026] = 642;
        test_data[2026] = 33'd2771483304;
        test_addr[2027] = 905;
        test_data[2027] = 33'd3962311491;
        test_addr[2028] = 944;
        test_data[2028] = 33'd4857802570;
        test_addr[2029] = 14;
        test_data[2029] = 33'd6781540609;
        test_addr[2030] = 140;
        test_data[2030] = 33'd8369234334;
        test_addr[2031] = 504;
        test_data[2031] = 33'd638967831;
        test_addr[2032] = 917;
        test_data[2032] = 33'd778607413;
        test_addr[2033] = 993;
        test_data[2033] = 33'd6873103799;
        test_addr[2034] = 815;
        test_data[2034] = 33'd4680758760;
        test_addr[2035] = 300;
        test_data[2035] = 33'd1695058610;
        test_addr[2036] = 483;
        test_data[2036] = 33'd4068064513;
        test_addr[2037] = 179;
        test_data[2037] = 33'd3882480974;
        test_addr[2038] = 595;
        test_data[2038] = 33'd2905081443;
        test_addr[2039] = 819;
        test_data[2039] = 33'd1860351677;
        test_addr[2040] = 933;
        test_data[2040] = 33'd4542305129;
        test_addr[2041] = 938;
        test_data[2041] = 33'd53485639;
        test_addr[2042] = 1006;
        test_data[2042] = 33'd904820223;
        test_addr[2043] = 968;
        test_data[2043] = 33'd3848370431;
        test_addr[2044] = 278;
        test_data[2044] = 33'd2148021305;
        test_addr[2045] = 638;
        test_data[2045] = 33'd5233924996;
        test_addr[2046] = 563;
        test_data[2046] = 33'd3249157073;
        test_addr[2047] = 921;
        test_data[2047] = 33'd7692955444;
        test_addr[2048] = 523;
        test_data[2048] = 33'd1209225517;
        test_addr[2049] = 488;
        test_data[2049] = 33'd1193364021;
        test_addr[2050] = 748;
        test_data[2050] = 33'd2905536779;
        test_addr[2051] = 294;
        test_data[2051] = 33'd301140059;
        test_addr[2052] = 257;
        test_data[2052] = 33'd4785507920;
        test_addr[2053] = 409;
        test_data[2053] = 33'd1379904639;
        test_addr[2054] = 923;
        test_data[2054] = 33'd412824823;
        test_addr[2055] = 620;
        test_data[2055] = 33'd990877164;
        test_addr[2056] = 267;
        test_data[2056] = 33'd904777788;
        test_addr[2057] = 387;
        test_data[2057] = 33'd2723287972;
        test_addr[2058] = 298;
        test_data[2058] = 33'd7701997189;
        test_addr[2059] = 144;
        test_data[2059] = 33'd3416637777;
        test_addr[2060] = 358;
        test_data[2060] = 33'd8467541585;
        test_addr[2061] = 358;
        test_data[2061] = 33'd4172574289;
        test_addr[2062] = 458;
        test_data[2062] = 33'd1978411341;
        test_addr[2063] = 888;
        test_data[2063] = 33'd4980958850;
        test_addr[2064] = 219;
        test_data[2064] = 33'd5218399040;
        test_addr[2065] = 359;
        test_data[2065] = 33'd3381025996;
        test_addr[2066] = 240;
        test_data[2066] = 33'd4066667004;
        test_addr[2067] = 18;
        test_data[2067] = 33'd4479556694;
        test_addr[2068] = 936;
        test_data[2068] = 33'd1292504590;
        test_addr[2069] = 262;
        test_data[2069] = 33'd8329244145;
        test_addr[2070] = 40;
        test_data[2070] = 33'd3594722951;
        test_addr[2071] = 4;
        test_data[2071] = 33'd1143739882;
        test_addr[2072] = 694;
        test_data[2072] = 33'd3417088654;
        test_addr[2073] = 960;
        test_data[2073] = 33'd5912451446;
        test_addr[2074] = 331;
        test_data[2074] = 33'd2402963099;
        test_addr[2075] = 478;
        test_data[2075] = 33'd2798923027;
        test_addr[2076] = 114;
        test_data[2076] = 33'd3622112771;
        test_addr[2077] = 991;
        test_data[2077] = 33'd1186657120;
        test_addr[2078] = 589;
        test_data[2078] = 33'd4364486303;
        test_addr[2079] = 967;
        test_data[2079] = 33'd8455836850;
        test_addr[2080] = 487;
        test_data[2080] = 33'd1196914595;
        test_addr[2081] = 573;
        test_data[2081] = 33'd3896166626;
        test_addr[2082] = 61;
        test_data[2082] = 33'd3050866392;
        test_addr[2083] = 824;
        test_data[2083] = 33'd403117584;
        test_addr[2084] = 490;
        test_data[2084] = 33'd1605742489;
        test_addr[2085] = 398;
        test_data[2085] = 33'd1613655084;
        test_addr[2086] = 732;
        test_data[2086] = 33'd1612454682;
        test_addr[2087] = 834;
        test_data[2087] = 33'd7085769886;
        test_addr[2088] = 705;
        test_data[2088] = 33'd3595301892;
        test_addr[2089] = 806;
        test_data[2089] = 33'd6875527619;
        test_addr[2090] = 1002;
        test_data[2090] = 33'd6654910697;
        test_addr[2091] = 646;
        test_data[2091] = 33'd132734761;
        test_addr[2092] = 938;
        test_data[2092] = 33'd53485639;
        test_addr[2093] = 228;
        test_data[2093] = 33'd1885599207;
        test_addr[2094] = 961;
        test_data[2094] = 33'd5761757774;
        test_addr[2095] = 952;
        test_data[2095] = 33'd6434304202;
        test_addr[2096] = 826;
        test_data[2096] = 33'd2881112742;
        test_addr[2097] = 580;
        test_data[2097] = 33'd4090953264;
        test_addr[2098] = 1013;
        test_data[2098] = 33'd3443847325;
        test_addr[2099] = 865;
        test_data[2099] = 33'd5965463068;
        test_addr[2100] = 602;
        test_data[2100] = 33'd5970007671;
        test_addr[2101] = 897;
        test_data[2101] = 33'd1039575909;
        test_addr[2102] = 948;
        test_data[2102] = 33'd3508169817;
        test_addr[2103] = 199;
        test_data[2103] = 33'd1949557997;
        test_addr[2104] = 700;
        test_data[2104] = 33'd2118661662;
        test_addr[2105] = 704;
        test_data[2105] = 33'd2828619334;
        test_addr[2106] = 976;
        test_data[2106] = 33'd3395753456;
        test_addr[2107] = 154;
        test_data[2107] = 33'd818530140;
        test_addr[2108] = 279;
        test_data[2108] = 33'd2094091315;
        test_addr[2109] = 575;
        test_data[2109] = 33'd4086039100;
        test_addr[2110] = 256;
        test_data[2110] = 33'd4365507330;
        test_addr[2111] = 448;
        test_data[2111] = 33'd2166151836;
        test_addr[2112] = 910;
        test_data[2112] = 33'd3948715188;
        test_addr[2113] = 333;
        test_data[2113] = 33'd3264659335;
        test_addr[2114] = 509;
        test_data[2114] = 33'd2005844869;
        test_addr[2115] = 191;
        test_data[2115] = 33'd3616306016;
        test_addr[2116] = 560;
        test_data[2116] = 33'd517678019;
        test_addr[2117] = 560;
        test_data[2117] = 33'd517678019;
        test_addr[2118] = 427;
        test_data[2118] = 33'd3283430231;
        test_addr[2119] = 455;
        test_data[2119] = 33'd4160999481;
        test_addr[2120] = 728;
        test_data[2120] = 33'd820874592;
        test_addr[2121] = 614;
        test_data[2121] = 33'd292281791;
        test_addr[2122] = 141;
        test_data[2122] = 33'd2186149626;
        test_addr[2123] = 187;
        test_data[2123] = 33'd1241473016;
        test_addr[2124] = 770;
        test_data[2124] = 33'd4502141641;
        test_addr[2125] = 8;
        test_data[2125] = 33'd3114571103;
        test_addr[2126] = 865;
        test_data[2126] = 33'd1670495772;
        test_addr[2127] = 730;
        test_data[2127] = 33'd7467152933;
        test_addr[2128] = 811;
        test_data[2128] = 33'd226245950;
        test_addr[2129] = 885;
        test_data[2129] = 33'd8360624052;
        test_addr[2130] = 634;
        test_data[2130] = 33'd5969177724;
        test_addr[2131] = 117;
        test_data[2131] = 33'd6723965449;
        test_addr[2132] = 731;
        test_data[2132] = 33'd914234311;
        test_addr[2133] = 717;
        test_data[2133] = 33'd2724895895;
        test_addr[2134] = 576;
        test_data[2134] = 33'd3521161878;
        test_addr[2135] = 1021;
        test_data[2135] = 33'd7158063905;
        test_addr[2136] = 614;
        test_data[2136] = 33'd5681611963;
        test_addr[2137] = 658;
        test_data[2137] = 33'd2510800920;
        test_addr[2138] = 682;
        test_data[2138] = 33'd3207157459;
        test_addr[2139] = 1010;
        test_data[2139] = 33'd6459089948;
        test_addr[2140] = 644;
        test_data[2140] = 33'd2060679594;
        test_addr[2141] = 991;
        test_data[2141] = 33'd1186657120;
        test_addr[2142] = 589;
        test_data[2142] = 33'd4949928888;
        test_addr[2143] = 189;
        test_data[2143] = 33'd5313695295;
        test_addr[2144] = 385;
        test_data[2144] = 33'd7032169256;
        test_addr[2145] = 831;
        test_data[2145] = 33'd2386706294;
        test_addr[2146] = 51;
        test_data[2146] = 33'd565760353;
        test_addr[2147] = 262;
        test_data[2147] = 33'd5345148894;
        test_addr[2148] = 303;
        test_data[2148] = 33'd3582560146;
        test_addr[2149] = 677;
        test_data[2149] = 33'd7091243556;
        test_addr[2150] = 130;
        test_data[2150] = 33'd939881898;
        test_addr[2151] = 86;
        test_data[2151] = 33'd2748145392;
        test_addr[2152] = 891;
        test_data[2152] = 33'd1858193830;
        test_addr[2153] = 41;
        test_data[2153] = 33'd786275004;
        test_addr[2154] = 29;
        test_data[2154] = 33'd1255285926;
        test_addr[2155] = 771;
        test_data[2155] = 33'd733190410;
        test_addr[2156] = 824;
        test_data[2156] = 33'd403117584;
        test_addr[2157] = 547;
        test_data[2157] = 33'd3532255610;
        test_addr[2158] = 841;
        test_data[2158] = 33'd8587004011;
        test_addr[2159] = 616;
        test_data[2159] = 33'd1933938369;
        test_addr[2160] = 732;
        test_data[2160] = 33'd5901743009;
        test_addr[2161] = 663;
        test_data[2161] = 33'd367404024;
        test_addr[2162] = 529;
        test_data[2162] = 33'd3797362521;
        test_addr[2163] = 356;
        test_data[2163] = 33'd6375652650;
        test_addr[2164] = 219;
        test_data[2164] = 33'd923431744;
        test_addr[2165] = 736;
        test_data[2165] = 33'd4060815809;
        test_addr[2166] = 122;
        test_data[2166] = 33'd5464498566;
        test_addr[2167] = 558;
        test_data[2167] = 33'd1054185022;
        test_addr[2168] = 373;
        test_data[2168] = 33'd8387230365;
        test_addr[2169] = 652;
        test_data[2169] = 33'd3345196147;
        test_addr[2170] = 974;
        test_data[2170] = 33'd3479926711;
        test_addr[2171] = 274;
        test_data[2171] = 33'd3059293611;
        test_addr[2172] = 378;
        test_data[2172] = 33'd1591577112;
        test_addr[2173] = 947;
        test_data[2173] = 33'd7216979296;
        test_addr[2174] = 816;
        test_data[2174] = 33'd2846493614;
        test_addr[2175] = 715;
        test_data[2175] = 33'd4108725227;
        test_addr[2176] = 101;
        test_data[2176] = 33'd334015143;
        test_addr[2177] = 926;
        test_data[2177] = 33'd4731000941;
        test_addr[2178] = 47;
        test_data[2178] = 33'd889566222;
        test_addr[2179] = 683;
        test_data[2179] = 33'd7078793614;
        test_addr[2180] = 82;
        test_data[2180] = 33'd2006336925;
        test_addr[2181] = 746;
        test_data[2181] = 33'd7962389891;
        test_addr[2182] = 680;
        test_data[2182] = 33'd1918095265;
        test_addr[2183] = 483;
        test_data[2183] = 33'd6646182813;
        test_addr[2184] = 157;
        test_data[2184] = 33'd5624102934;
        test_addr[2185] = 976;
        test_data[2185] = 33'd3395753456;
        test_addr[2186] = 55;
        test_data[2186] = 33'd812389879;
        test_addr[2187] = 51;
        test_data[2187] = 33'd565760353;
        test_addr[2188] = 965;
        test_data[2188] = 33'd8394343266;
        test_addr[2189] = 0;
        test_data[2189] = 33'd3077293961;
        test_addr[2190] = 529;
        test_data[2190] = 33'd3797362521;
        test_addr[2191] = 809;
        test_data[2191] = 33'd410675938;
        test_addr[2192] = 783;
        test_data[2192] = 33'd1379073191;
        test_addr[2193] = 383;
        test_data[2193] = 33'd1615749578;
        test_addr[2194] = 489;
        test_data[2194] = 33'd4219814471;
        test_addr[2195] = 301;
        test_data[2195] = 33'd3675695667;
        test_addr[2196] = 817;
        test_data[2196] = 33'd3133004597;
        test_addr[2197] = 302;
        test_data[2197] = 33'd1095590284;
        test_addr[2198] = 478;
        test_data[2198] = 33'd8168151309;
        test_addr[2199] = 691;
        test_data[2199] = 33'd3704402127;
        test_addr[2200] = 637;
        test_data[2200] = 33'd2030896509;
        test_addr[2201] = 881;
        test_data[2201] = 33'd2170563371;
        test_addr[2202] = 522;
        test_data[2202] = 33'd2055100449;
        test_addr[2203] = 725;
        test_data[2203] = 33'd4517436802;
        test_addr[2204] = 148;
        test_data[2204] = 33'd310279149;
        test_addr[2205] = 283;
        test_data[2205] = 33'd3321912760;
        test_addr[2206] = 311;
        test_data[2206] = 33'd1351719823;
        test_addr[2207] = 502;
        test_data[2207] = 33'd1213399919;
        test_addr[2208] = 709;
        test_data[2208] = 33'd2093977733;
        test_addr[2209] = 612;
        test_data[2209] = 33'd1343092192;
        test_addr[2210] = 908;
        test_data[2210] = 33'd3093603502;
        test_addr[2211] = 384;
        test_data[2211] = 33'd547271751;
        test_addr[2212] = 112;
        test_data[2212] = 33'd1757482678;
        test_addr[2213] = 295;
        test_data[2213] = 33'd2109502904;
        test_addr[2214] = 127;
        test_data[2214] = 33'd5561467461;
        test_addr[2215] = 84;
        test_data[2215] = 33'd5771901424;
        test_addr[2216] = 715;
        test_data[2216] = 33'd4108725227;
        test_addr[2217] = 334;
        test_data[2217] = 33'd4019955731;
        test_addr[2218] = 754;
        test_data[2218] = 33'd7073723442;
        test_addr[2219] = 766;
        test_data[2219] = 33'd1164223531;
        test_addr[2220] = 645;
        test_data[2220] = 33'd1478607793;
        test_addr[2221] = 786;
        test_data[2221] = 33'd4891706853;
        test_addr[2222] = 244;
        test_data[2222] = 33'd6825161738;
        test_addr[2223] = 715;
        test_data[2223] = 33'd6494304974;
        test_addr[2224] = 933;
        test_data[2224] = 33'd7333178268;
        test_addr[2225] = 809;
        test_data[2225] = 33'd7088751446;
        test_addr[2226] = 171;
        test_data[2226] = 33'd4662621770;
        test_addr[2227] = 870;
        test_data[2227] = 33'd8485135270;
        test_addr[2228] = 811;
        test_data[2228] = 33'd6653635035;
        test_addr[2229] = 368;
        test_data[2229] = 33'd329657286;
        test_addr[2230] = 733;
        test_data[2230] = 33'd1395512612;
        test_addr[2231] = 849;
        test_data[2231] = 33'd2242143770;
        test_addr[2232] = 356;
        test_data[2232] = 33'd7125367310;
        test_addr[2233] = 508;
        test_data[2233] = 33'd2458412144;
        test_addr[2234] = 350;
        test_data[2234] = 33'd2533041713;
        test_addr[2235] = 30;
        test_data[2235] = 33'd561337608;
        test_addr[2236] = 910;
        test_data[2236] = 33'd6128813262;
        test_addr[2237] = 743;
        test_data[2237] = 33'd6312086161;
        test_addr[2238] = 708;
        test_data[2238] = 33'd4183077687;
        test_addr[2239] = 851;
        test_data[2239] = 33'd1149027704;
        test_addr[2240] = 441;
        test_data[2240] = 33'd7902853733;
        test_addr[2241] = 162;
        test_data[2241] = 33'd1724568248;
        test_addr[2242] = 437;
        test_data[2242] = 33'd4732278737;
        test_addr[2243] = 860;
        test_data[2243] = 33'd562766076;
        test_addr[2244] = 307;
        test_data[2244] = 33'd6910169838;
        test_addr[2245] = 268;
        test_data[2245] = 33'd7187985233;
        test_addr[2246] = 398;
        test_data[2246] = 33'd5096176547;
        test_addr[2247] = 637;
        test_data[2247] = 33'd8340861975;
        test_addr[2248] = 103;
        test_data[2248] = 33'd3519285150;
        test_addr[2249] = 809;
        test_data[2249] = 33'd2793784150;
        test_addr[2250] = 257;
        test_data[2250] = 33'd490540624;
        test_addr[2251] = 154;
        test_data[2251] = 33'd818530140;
        test_addr[2252] = 1000;
        test_data[2252] = 33'd8187111692;
        test_addr[2253] = 862;
        test_data[2253] = 33'd1299278838;
        test_addr[2254] = 430;
        test_data[2254] = 33'd8144134942;
        test_addr[2255] = 938;
        test_data[2255] = 33'd53485639;
        test_addr[2256] = 903;
        test_data[2256] = 33'd3268229861;
        test_addr[2257] = 315;
        test_data[2257] = 33'd1859419918;
        test_addr[2258] = 881;
        test_data[2258] = 33'd2170563371;
        test_addr[2259] = 680;
        test_data[2259] = 33'd6295441502;
        test_addr[2260] = 437;
        test_data[2260] = 33'd437311441;
        test_addr[2261] = 322;
        test_data[2261] = 33'd26007573;
        test_addr[2262] = 188;
        test_data[2262] = 33'd5998907101;
        test_addr[2263] = 540;
        test_data[2263] = 33'd3411388360;
        test_addr[2264] = 339;
        test_data[2264] = 33'd3510710878;
        test_addr[2265] = 64;
        test_data[2265] = 33'd1257723553;
        test_addr[2266] = 707;
        test_data[2266] = 33'd1855980571;
        test_addr[2267] = 213;
        test_data[2267] = 33'd8440615901;
        test_addr[2268] = 360;
        test_data[2268] = 33'd7918328992;
        test_addr[2269] = 337;
        test_data[2269] = 33'd3555484088;
        test_addr[2270] = 729;
        test_data[2270] = 33'd1893345796;
        test_addr[2271] = 568;
        test_data[2271] = 33'd3549289617;
        test_addr[2272] = 159;
        test_data[2272] = 33'd3848464431;
        test_addr[2273] = 164;
        test_data[2273] = 33'd448429293;
        test_addr[2274] = 945;
        test_data[2274] = 33'd6088310710;
        test_addr[2275] = 771;
        test_data[2275] = 33'd733190410;
        test_addr[2276] = 944;
        test_data[2276] = 33'd7420942445;
        test_addr[2277] = 3;
        test_data[2277] = 33'd2710397198;
        test_addr[2278] = 803;
        test_data[2278] = 33'd7944188427;
        test_addr[2279] = 666;
        test_data[2279] = 33'd1952473218;
        test_addr[2280] = 87;
        test_data[2280] = 33'd3390580480;
        test_addr[2281] = 939;
        test_data[2281] = 33'd3724952086;
        test_addr[2282] = 617;
        test_data[2282] = 33'd306081816;
        test_addr[2283] = 147;
        test_data[2283] = 33'd5766961294;
        test_addr[2284] = 231;
        test_data[2284] = 33'd2571519824;
        test_addr[2285] = 7;
        test_data[2285] = 33'd2323112615;
        test_addr[2286] = 781;
        test_data[2286] = 33'd1625107923;
        test_addr[2287] = 1004;
        test_data[2287] = 33'd1981183283;
        test_addr[2288] = 45;
        test_data[2288] = 33'd1127328015;
        test_addr[2289] = 127;
        test_data[2289] = 33'd7232492334;
        test_addr[2290] = 41;
        test_data[2290] = 33'd786275004;
        test_addr[2291] = 657;
        test_data[2291] = 33'd927834072;
        test_addr[2292] = 382;
        test_data[2292] = 33'd706838701;
        test_addr[2293] = 193;
        test_data[2293] = 33'd7887274045;
        test_addr[2294] = 696;
        test_data[2294] = 33'd7837075157;
        test_addr[2295] = 37;
        test_data[2295] = 33'd8504520160;
        test_addr[2296] = 12;
        test_data[2296] = 33'd1981417174;
        test_addr[2297] = 492;
        test_data[2297] = 33'd4265285582;
        test_addr[2298] = 35;
        test_data[2298] = 33'd3955127962;
        test_addr[2299] = 113;
        test_data[2299] = 33'd5364652406;
        test_addr[2300] = 1005;
        test_data[2300] = 33'd3281370832;
        test_addr[2301] = 1002;
        test_data[2301] = 33'd2359943401;
        test_addr[2302] = 470;
        test_data[2302] = 33'd4198953116;
        test_addr[2303] = 721;
        test_data[2303] = 33'd3714234635;
        test_addr[2304] = 82;
        test_data[2304] = 33'd2006336925;
        test_addr[2305] = 821;
        test_data[2305] = 33'd2331168722;
        test_addr[2306] = 475;
        test_data[2306] = 33'd2559009820;
        test_addr[2307] = 162;
        test_data[2307] = 33'd1724568248;
        test_addr[2308] = 293;
        test_data[2308] = 33'd2329958859;
        test_addr[2309] = 354;
        test_data[2309] = 33'd1554725479;
        test_addr[2310] = 504;
        test_data[2310] = 33'd638967831;
        test_addr[2311] = 561;
        test_data[2311] = 33'd7392603853;
        test_addr[2312] = 14;
        test_data[2312] = 33'd2486573313;
        test_addr[2313] = 913;
        test_data[2313] = 33'd5098256723;
        test_addr[2314] = 425;
        test_data[2314] = 33'd3413574269;
        test_addr[2315] = 11;
        test_data[2315] = 33'd1048550729;
        test_addr[2316] = 815;
        test_data[2316] = 33'd385791464;
        test_addr[2317] = 524;
        test_data[2317] = 33'd527412138;
        test_addr[2318] = 812;
        test_data[2318] = 33'd2158247624;
        test_addr[2319] = 832;
        test_data[2319] = 33'd4621416576;
        test_addr[2320] = 174;
        test_data[2320] = 33'd5159150941;
        test_addr[2321] = 848;
        test_data[2321] = 33'd74868948;
        test_addr[2322] = 896;
        test_data[2322] = 33'd3066857618;
        test_addr[2323] = 692;
        test_data[2323] = 33'd8214207815;
        test_addr[2324] = 591;
        test_data[2324] = 33'd6849075480;
        test_addr[2325] = 540;
        test_data[2325] = 33'd8125214370;
        test_addr[2326] = 117;
        test_data[2326] = 33'd2428998153;
        test_addr[2327] = 758;
        test_data[2327] = 33'd1957858034;
        test_addr[2328] = 786;
        test_data[2328] = 33'd596739557;
        test_addr[2329] = 86;
        test_data[2329] = 33'd2748145392;
        test_addr[2330] = 883;
        test_data[2330] = 33'd43240007;
        test_addr[2331] = 722;
        test_data[2331] = 33'd6957426088;
        test_addr[2332] = 256;
        test_data[2332] = 33'd5140603855;
        test_addr[2333] = 215;
        test_data[2333] = 33'd815101909;
        test_addr[2334] = 825;
        test_data[2334] = 33'd4252998212;
        test_addr[2335] = 938;
        test_data[2335] = 33'd6529453995;
        test_addr[2336] = 498;
        test_data[2336] = 33'd3710558399;
        test_addr[2337] = 429;
        test_data[2337] = 33'd5696598689;
        test_addr[2338] = 270;
        test_data[2338] = 33'd8587214499;
        test_addr[2339] = 929;
        test_data[2339] = 33'd2524469636;
        test_addr[2340] = 562;
        test_data[2340] = 33'd4854839457;
        test_addr[2341] = 912;
        test_data[2341] = 33'd1730083639;
        test_addr[2342] = 483;
        test_data[2342] = 33'd5237895541;
        test_addr[2343] = 295;
        test_data[2343] = 33'd2109502904;
        test_addr[2344] = 830;
        test_data[2344] = 33'd3539273762;
        test_addr[2345] = 380;
        test_data[2345] = 33'd2260081304;
        test_addr[2346] = 636;
        test_data[2346] = 33'd1854299730;
        test_addr[2347] = 286;
        test_data[2347] = 33'd5478511028;
        test_addr[2348] = 78;
        test_data[2348] = 33'd3865815998;
        test_addr[2349] = 695;
        test_data[2349] = 33'd1994408553;
        test_addr[2350] = 913;
        test_data[2350] = 33'd803289427;
        test_addr[2351] = 939;
        test_data[2351] = 33'd3724952086;
        test_addr[2352] = 869;
        test_data[2352] = 33'd7873526532;
        test_addr[2353] = 204;
        test_data[2353] = 33'd2557857253;
        test_addr[2354] = 520;
        test_data[2354] = 33'd2224233289;
        test_addr[2355] = 589;
        test_data[2355] = 33'd654961592;
        test_addr[2356] = 366;
        test_data[2356] = 33'd2558372418;
        test_addr[2357] = 666;
        test_data[2357] = 33'd1952473218;
        test_addr[2358] = 279;
        test_data[2358] = 33'd2094091315;
        test_addr[2359] = 742;
        test_data[2359] = 33'd5472074167;
        test_addr[2360] = 647;
        test_data[2360] = 33'd1466466644;
        test_addr[2361] = 185;
        test_data[2361] = 33'd3678596044;
        test_addr[2362] = 975;
        test_data[2362] = 33'd4004751704;
        test_addr[2363] = 189;
        test_data[2363] = 33'd5128360337;
        test_addr[2364] = 951;
        test_data[2364] = 33'd2460043506;
        test_addr[2365] = 472;
        test_data[2365] = 33'd794664940;
        test_addr[2366] = 331;
        test_data[2366] = 33'd2402963099;
        test_addr[2367] = 850;
        test_data[2367] = 33'd2610616633;
        test_addr[2368] = 947;
        test_data[2368] = 33'd2922012000;
        test_addr[2369] = 895;
        test_data[2369] = 33'd7383934296;
        test_addr[2370] = 902;
        test_data[2370] = 33'd1242100171;
        test_addr[2371] = 775;
        test_data[2371] = 33'd1688794719;
        test_addr[2372] = 817;
        test_data[2372] = 33'd3133004597;
        test_addr[2373] = 317;
        test_data[2373] = 33'd2142036855;
        test_addr[2374] = 512;
        test_data[2374] = 33'd4210439056;
        test_addr[2375] = 669;
        test_data[2375] = 33'd459165770;
        test_addr[2376] = 93;
        test_data[2376] = 33'd3012159401;
        test_addr[2377] = 782;
        test_data[2377] = 33'd2982764277;
        test_addr[2378] = 197;
        test_data[2378] = 33'd4143794548;
        test_addr[2379] = 60;
        test_data[2379] = 33'd1436918879;
        test_addr[2380] = 410;
        test_data[2380] = 33'd3670908267;
        test_addr[2381] = 1006;
        test_data[2381] = 33'd904820223;
        test_addr[2382] = 453;
        test_data[2382] = 33'd3500901833;
        test_addr[2383] = 18;
        test_data[2383] = 33'd7315295882;
        test_addr[2384] = 23;
        test_data[2384] = 33'd2328303965;
        test_addr[2385] = 131;
        test_data[2385] = 33'd3754095223;
        test_addr[2386] = 354;
        test_data[2386] = 33'd1554725479;
        test_addr[2387] = 31;
        test_data[2387] = 33'd2160288399;
        test_addr[2388] = 377;
        test_data[2388] = 33'd7448110148;
        test_addr[2389] = 558;
        test_data[2389] = 33'd1054185022;
        test_addr[2390] = 975;
        test_data[2390] = 33'd5416575199;
        test_addr[2391] = 90;
        test_data[2391] = 33'd684440951;
        test_addr[2392] = 624;
        test_data[2392] = 33'd2766751231;
        test_addr[2393] = 682;
        test_data[2393] = 33'd3207157459;
        test_addr[2394] = 60;
        test_data[2394] = 33'd6587968892;
        test_addr[2395] = 612;
        test_data[2395] = 33'd5132783025;
        test_addr[2396] = 178;
        test_data[2396] = 33'd3708009236;
        test_addr[2397] = 589;
        test_data[2397] = 33'd654961592;
        test_addr[2398] = 11;
        test_data[2398] = 33'd6639302387;
        test_addr[2399] = 37;
        test_data[2399] = 33'd4209552864;
        test_addr[2400] = 140;
        test_data[2400] = 33'd4074267038;
        test_addr[2401] = 569;
        test_data[2401] = 33'd2633019442;
        test_addr[2402] = 569;
        test_data[2402] = 33'd2633019442;
        test_addr[2403] = 585;
        test_data[2403] = 33'd8368045370;
        test_addr[2404] = 957;
        test_data[2404] = 33'd4600050734;
        test_addr[2405] = 215;
        test_data[2405] = 33'd5322938906;
        test_addr[2406] = 587;
        test_data[2406] = 33'd3580683813;
        test_addr[2407] = 3;
        test_data[2407] = 33'd2710397198;
        test_addr[2408] = 636;
        test_data[2408] = 33'd1854299730;
        test_addr[2409] = 380;
        test_data[2409] = 33'd2260081304;
        test_addr[2410] = 488;
        test_data[2410] = 33'd1193364021;
        test_addr[2411] = 763;
        test_data[2411] = 33'd1119246121;
        test_addr[2412] = 549;
        test_data[2412] = 33'd3183535881;
        test_addr[2413] = 292;
        test_data[2413] = 33'd1265860839;
        test_addr[2414] = 828;
        test_data[2414] = 33'd1107521268;
        test_addr[2415] = 255;
        test_data[2415] = 33'd7191962577;
        test_addr[2416] = 414;
        test_data[2416] = 33'd7419845935;
        test_addr[2417] = 49;
        test_data[2417] = 33'd1117414700;
        test_addr[2418] = 267;
        test_data[2418] = 33'd904777788;
        test_addr[2419] = 2;
        test_data[2419] = 33'd2348039952;
        test_addr[2420] = 577;
        test_data[2420] = 33'd2874325634;
        test_addr[2421] = 30;
        test_data[2421] = 33'd561337608;
        test_addr[2422] = 397;
        test_data[2422] = 33'd4518768614;
        test_addr[2423] = 183;
        test_data[2423] = 33'd4442843;
        test_addr[2424] = 906;
        test_data[2424] = 33'd3294149566;
        test_addr[2425] = 774;
        test_data[2425] = 33'd5618238874;
        test_addr[2426] = 835;
        test_data[2426] = 33'd1686846772;
        test_addr[2427] = 59;
        test_data[2427] = 33'd1947913714;
        test_addr[2428] = 361;
        test_data[2428] = 33'd1290055053;
        test_addr[2429] = 925;
        test_data[2429] = 33'd1219013972;
        test_addr[2430] = 494;
        test_data[2430] = 33'd1860698751;
        test_addr[2431] = 245;
        test_data[2431] = 33'd1366539889;
        test_addr[2432] = 122;
        test_data[2432] = 33'd5782041101;
        test_addr[2433] = 856;
        test_data[2433] = 33'd2857576750;
        test_addr[2434] = 806;
        test_data[2434] = 33'd2580560323;
        test_addr[2435] = 357;
        test_data[2435] = 33'd2986504088;
        test_addr[2436] = 933;
        test_data[2436] = 33'd3038210972;
        test_addr[2437] = 353;
        test_data[2437] = 33'd1320710077;
        test_addr[2438] = 776;
        test_data[2438] = 33'd2409863467;
        test_addr[2439] = 344;
        test_data[2439] = 33'd6282016420;
        test_addr[2440] = 35;
        test_data[2440] = 33'd3955127962;
        test_addr[2441] = 494;
        test_data[2441] = 33'd1860698751;
        test_addr[2442] = 116;
        test_data[2442] = 33'd8211828913;
        test_addr[2443] = 317;
        test_data[2443] = 33'd2142036855;
        test_addr[2444] = 868;
        test_data[2444] = 33'd2145195459;
        test_addr[2445] = 602;
        test_data[2445] = 33'd1675040375;
        test_addr[2446] = 229;
        test_data[2446] = 33'd1480893710;
        test_addr[2447] = 228;
        test_data[2447] = 33'd1885599207;
        test_addr[2448] = 86;
        test_data[2448] = 33'd5431052556;
        test_addr[2449] = 844;
        test_data[2449] = 33'd6280780172;
        test_addr[2450] = 525;
        test_data[2450] = 33'd3648823425;
        test_addr[2451] = 219;
        test_data[2451] = 33'd923431744;
        test_addr[2452] = 458;
        test_data[2452] = 33'd1978411341;
        test_addr[2453] = 773;
        test_data[2453] = 33'd531933772;
        test_addr[2454] = 115;
        test_data[2454] = 33'd4938645312;
        test_addr[2455] = 313;
        test_data[2455] = 33'd2220400995;
        test_addr[2456] = 549;
        test_data[2456] = 33'd3183535881;
        test_addr[2457] = 101;
        test_data[2457] = 33'd334015143;
        test_addr[2458] = 492;
        test_data[2458] = 33'd4265285582;
        test_addr[2459] = 293;
        test_data[2459] = 33'd2329958859;
        test_addr[2460] = 508;
        test_data[2460] = 33'd8095388447;
        test_addr[2461] = 49;
        test_data[2461] = 33'd5590513085;
        test_addr[2462] = 641;
        test_data[2462] = 33'd6531508555;
        test_addr[2463] = 354;
        test_data[2463] = 33'd1554725479;
        test_addr[2464] = 193;
        test_data[2464] = 33'd5381752294;
        test_addr[2465] = 758;
        test_data[2465] = 33'd1957858034;
        test_addr[2466] = 208;
        test_data[2466] = 33'd881023582;
        test_addr[2467] = 153;
        test_data[2467] = 33'd1670173968;
        test_addr[2468] = 38;
        test_data[2468] = 33'd1762764931;
        test_addr[2469] = 498;
        test_data[2469] = 33'd5612860127;
        test_addr[2470] = 227;
        test_data[2470] = 33'd8409021968;
        test_addr[2471] = 864;
        test_data[2471] = 33'd702666674;
        test_addr[2472] = 363;
        test_data[2472] = 33'd3448701357;
        test_addr[2473] = 969;
        test_data[2473] = 33'd1593693352;
        test_addr[2474] = 125;
        test_data[2474] = 33'd5554701001;
        test_addr[2475] = 44;
        test_data[2475] = 33'd3885394360;
        test_addr[2476] = 812;
        test_data[2476] = 33'd2158247624;
        test_addr[2477] = 886;
        test_data[2477] = 33'd479387173;
        test_addr[2478] = 300;
        test_data[2478] = 33'd6815243567;
        test_addr[2479] = 335;
        test_data[2479] = 33'd7692253651;
        test_addr[2480] = 145;
        test_data[2480] = 33'd200240380;
        test_addr[2481] = 623;
        test_data[2481] = 33'd4276947268;
        test_addr[2482] = 656;
        test_data[2482] = 33'd4186206039;
        test_addr[2483] = 866;
        test_data[2483] = 33'd2619727747;
        test_addr[2484] = 242;
        test_data[2484] = 33'd2171707476;
        test_addr[2485] = 384;
        test_data[2485] = 33'd547271751;
        test_addr[2486] = 1020;
        test_data[2486] = 33'd3144327154;
        test_addr[2487] = 541;
        test_data[2487] = 33'd2903716974;
        test_addr[2488] = 173;
        test_data[2488] = 33'd4580647132;
        test_addr[2489] = 485;
        test_data[2489] = 33'd4058835011;
        test_addr[2490] = 573;
        test_data[2490] = 33'd3896166626;
        test_addr[2491] = 705;
        test_data[2491] = 33'd5392524722;
        test_addr[2492] = 540;
        test_data[2492] = 33'd3830247074;
        test_addr[2493] = 579;
        test_data[2493] = 33'd7245534812;
        test_addr[2494] = 394;
        test_data[2494] = 33'd2134209481;
        test_addr[2495] = 896;
        test_data[2495] = 33'd7917824911;
        test_addr[2496] = 670;
        test_data[2496] = 33'd7700420448;
        test_addr[2497] = 285;
        test_data[2497] = 33'd6138026938;
        test_addr[2498] = 787;
        test_data[2498] = 33'd2332338642;
        test_addr[2499] = 480;
        test_data[2499] = 33'd2118543923;
        test_addr[2500] = 747;
        test_data[2500] = 33'd901675206;
        test_addr[2501] = 349;
        test_data[2501] = 33'd394458336;
        test_addr[2502] = 534;
        test_data[2502] = 33'd3992358006;
        test_addr[2503] = 847;
        test_data[2503] = 33'd1925753163;
        test_addr[2504] = 322;
        test_data[2504] = 33'd26007573;
        test_addr[2505] = 979;
        test_data[2505] = 33'd4522222612;
        test_addr[2506] = 963;
        test_data[2506] = 33'd4567587591;
        test_addr[2507] = 185;
        test_data[2507] = 33'd5099566863;
        test_addr[2508] = 837;
        test_data[2508] = 33'd1693487156;
        test_addr[2509] = 39;
        test_data[2509] = 33'd5957107320;
        test_addr[2510] = 799;
        test_data[2510] = 33'd4497021828;
        test_addr[2511] = 61;
        test_data[2511] = 33'd3050866392;
        test_addr[2512] = 870;
        test_data[2512] = 33'd5543970508;
        test_addr[2513] = 899;
        test_data[2513] = 33'd5356371113;
        test_addr[2514] = 793;
        test_data[2514] = 33'd5157853656;
        test_addr[2515] = 187;
        test_data[2515] = 33'd6905827359;
        test_addr[2516] = 74;
        test_data[2516] = 33'd5892408442;
        test_addr[2517] = 51;
        test_data[2517] = 33'd565760353;
        test_addr[2518] = 59;
        test_data[2518] = 33'd1947913714;
        test_addr[2519] = 350;
        test_data[2519] = 33'd2533041713;
        test_addr[2520] = 319;
        test_data[2520] = 33'd3354761559;
        test_addr[2521] = 50;
        test_data[2521] = 33'd1824887721;
        test_addr[2522] = 308;
        test_data[2522] = 33'd2304201728;
        test_addr[2523] = 666;
        test_data[2523] = 33'd7737514309;
        test_addr[2524] = 679;
        test_data[2524] = 33'd2110703835;
        test_addr[2525] = 554;
        test_data[2525] = 33'd4310766579;
        test_addr[2526] = 586;
        test_data[2526] = 33'd5898570520;
        test_addr[2527] = 293;
        test_data[2527] = 33'd2329958859;
        test_addr[2528] = 813;
        test_data[2528] = 33'd5903376117;
        test_addr[2529] = 289;
        test_data[2529] = 33'd3920997515;
        test_addr[2530] = 239;
        test_data[2530] = 33'd4506925806;
        test_addr[2531] = 370;
        test_data[2531] = 33'd4079085858;
        test_addr[2532] = 835;
        test_data[2532] = 33'd4430813258;
        test_addr[2533] = 414;
        test_data[2533] = 33'd7866184270;
        test_addr[2534] = 891;
        test_data[2534] = 33'd1858193830;
        test_addr[2535] = 636;
        test_data[2535] = 33'd1854299730;
        test_addr[2536] = 415;
        test_data[2536] = 33'd95744961;
        test_addr[2537] = 795;
        test_data[2537] = 33'd88944858;
        test_addr[2538] = 37;
        test_data[2538] = 33'd4328547467;
        test_addr[2539] = 555;
        test_data[2539] = 33'd1371209800;
        test_addr[2540] = 265;
        test_data[2540] = 33'd6100436917;
        test_addr[2541] = 612;
        test_data[2541] = 33'd837815729;
        test_addr[2542] = 765;
        test_data[2542] = 33'd843852261;
        test_addr[2543] = 386;
        test_data[2543] = 33'd7596117821;
        test_addr[2544] = 345;
        test_data[2544] = 33'd8067540263;
        test_addr[2545] = 68;
        test_data[2545] = 33'd780007243;
        test_addr[2546] = 662;
        test_data[2546] = 33'd4544273189;
        test_addr[2547] = 686;
        test_data[2547] = 33'd4286094390;
        test_addr[2548] = 446;
        test_data[2548] = 33'd1055605986;
        test_addr[2549] = 638;
        test_data[2549] = 33'd938957700;
        test_addr[2550] = 109;
        test_data[2550] = 33'd2687315092;
        test_addr[2551] = 262;
        test_data[2551] = 33'd1050181598;
        test_addr[2552] = 739;
        test_data[2552] = 33'd24113143;
        test_addr[2553] = 1023;
        test_data[2553] = 33'd107160650;
        test_addr[2554] = 239;
        test_data[2554] = 33'd7603507020;
        test_addr[2555] = 276;
        test_data[2555] = 33'd1049188557;
        test_addr[2556] = 157;
        test_data[2556] = 33'd5205809401;
        test_addr[2557] = 836;
        test_data[2557] = 33'd4656346490;
        test_addr[2558] = 477;
        test_data[2558] = 33'd4727966373;
        test_addr[2559] = 168;
        test_data[2559] = 33'd6951801890;
        test_addr[2560] = 829;
        test_data[2560] = 33'd7046161648;
        test_addr[2561] = 743;
        test_data[2561] = 33'd5034013001;
        test_addr[2562] = 728;
        test_data[2562] = 33'd6665371184;
        test_addr[2563] = 79;
        test_data[2563] = 33'd4243798425;
        test_addr[2564] = 731;
        test_data[2564] = 33'd4647688567;
        test_addr[2565] = 202;
        test_data[2565] = 33'd2314598239;
        test_addr[2566] = 798;
        test_data[2566] = 33'd4210928188;
        test_addr[2567] = 149;
        test_data[2567] = 33'd96483764;
        test_addr[2568] = 7;
        test_data[2568] = 33'd5352983526;
        test_addr[2569] = 765;
        test_data[2569] = 33'd843852261;
        test_addr[2570] = 496;
        test_data[2570] = 33'd262877978;
        test_addr[2571] = 414;
        test_data[2571] = 33'd7888561034;
        test_addr[2572] = 491;
        test_data[2572] = 33'd6033685137;
        test_addr[2573] = 576;
        test_data[2573] = 33'd3521161878;
        test_addr[2574] = 35;
        test_data[2574] = 33'd3955127962;
        test_addr[2575] = 206;
        test_data[2575] = 33'd3440932254;
        test_addr[2576] = 428;
        test_data[2576] = 33'd192890954;
        test_addr[2577] = 803;
        test_data[2577] = 33'd4397431513;
        test_addr[2578] = 565;
        test_data[2578] = 33'd4241384530;
        test_addr[2579] = 103;
        test_data[2579] = 33'd8385607166;
        test_addr[2580] = 502;
        test_data[2580] = 33'd1213399919;
        test_addr[2581] = 872;
        test_data[2581] = 33'd8000286110;
        test_addr[2582] = 876;
        test_data[2582] = 33'd1222913046;
        test_addr[2583] = 743;
        test_data[2583] = 33'd739045705;
        test_addr[2584] = 765;
        test_data[2584] = 33'd843852261;
        test_addr[2585] = 369;
        test_data[2585] = 33'd3108046467;
        test_addr[2586] = 265;
        test_data[2586] = 33'd1805469621;
        test_addr[2587] = 47;
        test_data[2587] = 33'd889566222;
        test_addr[2588] = 945;
        test_data[2588] = 33'd1793343414;
        test_addr[2589] = 882;
        test_data[2589] = 33'd2715226243;
        test_addr[2590] = 281;
        test_data[2590] = 33'd8403670296;
        test_addr[2591] = 309;
        test_data[2591] = 33'd2815024490;
        test_addr[2592] = 821;
        test_data[2592] = 33'd7450995738;
        test_addr[2593] = 926;
        test_data[2593] = 33'd436033645;
        test_addr[2594] = 22;
        test_data[2594] = 33'd2308919392;
        test_addr[2595] = 809;
        test_data[2595] = 33'd4524560550;
        test_addr[2596] = 936;
        test_data[2596] = 33'd1292504590;
        test_addr[2597] = 515;
        test_data[2597] = 33'd183309785;
        test_addr[2598] = 974;
        test_data[2598] = 33'd3479926711;
        test_addr[2599] = 967;
        test_data[2599] = 33'd4160869554;
        test_addr[2600] = 69;
        test_data[2600] = 33'd5970217936;
        test_addr[2601] = 131;
        test_data[2601] = 33'd3754095223;
        test_addr[2602] = 1010;
        test_data[2602] = 33'd2164122652;
        test_addr[2603] = 851;
        test_data[2603] = 33'd5147093866;
        test_addr[2604] = 158;
        test_data[2604] = 33'd370641019;
        test_addr[2605] = 654;
        test_data[2605] = 33'd984783600;
        test_addr[2606] = 797;
        test_data[2606] = 33'd3094034019;
        test_addr[2607] = 627;
        test_data[2607] = 33'd2656035837;
        test_addr[2608] = 769;
        test_data[2608] = 33'd3111199946;
        test_addr[2609] = 206;
        test_data[2609] = 33'd3440932254;
        test_addr[2610] = 161;
        test_data[2610] = 33'd1596641998;
        test_addr[2611] = 517;
        test_data[2611] = 33'd441152082;
        test_addr[2612] = 371;
        test_data[2612] = 33'd768853880;
        test_addr[2613] = 975;
        test_data[2613] = 33'd8546851599;
        test_addr[2614] = 700;
        test_data[2614] = 33'd2118661662;
        test_addr[2615] = 978;
        test_data[2615] = 33'd1849704765;
        test_addr[2616] = 645;
        test_data[2616] = 33'd4538838748;
        test_addr[2617] = 622;
        test_data[2617] = 33'd3997591646;
        test_addr[2618] = 571;
        test_data[2618] = 33'd6849695852;
        test_addr[2619] = 872;
        test_data[2619] = 33'd3705318814;
        test_addr[2620] = 509;
        test_data[2620] = 33'd2005844869;
        test_addr[2621] = 251;
        test_data[2621] = 33'd3084835230;
        test_addr[2622] = 597;
        test_data[2622] = 33'd2521741564;
        test_addr[2623] = 512;
        test_data[2623] = 33'd4210439056;
        test_addr[2624] = 186;
        test_data[2624] = 33'd4050893006;
        test_addr[2625] = 719;
        test_data[2625] = 33'd6971209281;
        test_addr[2626] = 684;
        test_data[2626] = 33'd300267709;
        test_addr[2627] = 114;
        test_data[2627] = 33'd3622112771;
        test_addr[2628] = 449;
        test_data[2628] = 33'd6693894183;
        test_addr[2629] = 94;
        test_data[2629] = 33'd549339061;
        test_addr[2630] = 242;
        test_data[2630] = 33'd2171707476;
        test_addr[2631] = 105;
        test_data[2631] = 33'd1192418195;
        test_addr[2632] = 746;
        test_data[2632] = 33'd3667422595;
        test_addr[2633] = 1019;
        test_data[2633] = 33'd510091675;
        test_addr[2634] = 144;
        test_data[2634] = 33'd3416637777;
        test_addr[2635] = 867;
        test_data[2635] = 33'd1994039453;
        test_addr[2636] = 789;
        test_data[2636] = 33'd5251398752;
        test_addr[2637] = 24;
        test_data[2637] = 33'd5972863267;
        test_addr[2638] = 983;
        test_data[2638] = 33'd8326877364;
        test_addr[2639] = 431;
        test_data[2639] = 33'd2717572314;
        test_addr[2640] = 391;
        test_data[2640] = 33'd3059314876;
        test_addr[2641] = 638;
        test_data[2641] = 33'd5462636952;
        test_addr[2642] = 225;
        test_data[2642] = 33'd524980437;
        test_addr[2643] = 1003;
        test_data[2643] = 33'd6962279107;
        test_addr[2644] = 990;
        test_data[2644] = 33'd616895957;
        test_addr[2645] = 652;
        test_data[2645] = 33'd3345196147;
        test_addr[2646] = 846;
        test_data[2646] = 33'd258233883;
        test_addr[2647] = 662;
        test_data[2647] = 33'd249305893;
        test_addr[2648] = 141;
        test_data[2648] = 33'd2186149626;
        test_addr[2649] = 369;
        test_data[2649] = 33'd5819687681;
        test_addr[2650] = 1015;
        test_data[2650] = 33'd8228804880;
        test_addr[2651] = 667;
        test_data[2651] = 33'd7738714675;
        test_addr[2652] = 205;
        test_data[2652] = 33'd8334869082;
        test_addr[2653] = 811;
        test_data[2653] = 33'd2358667739;
        test_addr[2654] = 503;
        test_data[2654] = 33'd3936231662;
        test_addr[2655] = 49;
        test_data[2655] = 33'd8496863574;
        test_addr[2656] = 355;
        test_data[2656] = 33'd6886475090;
        test_addr[2657] = 624;
        test_data[2657] = 33'd2766751231;
        test_addr[2658] = 678;
        test_data[2658] = 33'd3688685586;
        test_addr[2659] = 149;
        test_data[2659] = 33'd96483764;
        test_addr[2660] = 191;
        test_data[2660] = 33'd3616306016;
        test_addr[2661] = 233;
        test_data[2661] = 33'd1331185298;
        test_addr[2662] = 640;
        test_data[2662] = 33'd7275105657;
        test_addr[2663] = 487;
        test_data[2663] = 33'd4571088211;
        test_addr[2664] = 76;
        test_data[2664] = 33'd648789103;
        test_addr[2665] = 128;
        test_data[2665] = 33'd2369463817;
        test_addr[2666] = 573;
        test_data[2666] = 33'd3896166626;
        test_addr[2667] = 368;
        test_data[2667] = 33'd329657286;
        test_addr[2668] = 461;
        test_data[2668] = 33'd8089064603;
        test_addr[2669] = 822;
        test_data[2669] = 33'd3946742381;
        test_addr[2670] = 375;
        test_data[2670] = 33'd5091936292;
        test_addr[2671] = 59;
        test_data[2671] = 33'd1947913714;
        test_addr[2672] = 84;
        test_data[2672] = 33'd1476934128;
        test_addr[2673] = 58;
        test_data[2673] = 33'd2543580284;
        test_addr[2674] = 172;
        test_data[2674] = 33'd3528050181;
        test_addr[2675] = 823;
        test_data[2675] = 33'd700710660;
        test_addr[2676] = 983;
        test_data[2676] = 33'd4031910068;
        test_addr[2677] = 947;
        test_data[2677] = 33'd2922012000;
        test_addr[2678] = 930;
        test_data[2678] = 33'd5658964965;
        test_addr[2679] = 747;
        test_data[2679] = 33'd901675206;
        test_addr[2680] = 1009;
        test_data[2680] = 33'd3939855400;
        test_addr[2681] = 674;
        test_data[2681] = 33'd1833629200;
        test_addr[2682] = 379;
        test_data[2682] = 33'd7504310587;
        test_addr[2683] = 374;
        test_data[2683] = 33'd2803425201;
        test_addr[2684] = 758;
        test_data[2684] = 33'd7652110259;
        test_addr[2685] = 930;
        test_data[2685] = 33'd1363997669;
        test_addr[2686] = 286;
        test_data[2686] = 33'd6576952045;
        test_addr[2687] = 69;
        test_data[2687] = 33'd1675250640;
        test_addr[2688] = 744;
        test_data[2688] = 33'd2105270382;
        test_addr[2689] = 14;
        test_data[2689] = 33'd2486573313;
        test_addr[2690] = 473;
        test_data[2690] = 33'd2897863862;
        test_addr[2691] = 501;
        test_data[2691] = 33'd138578467;
        test_addr[2692] = 266;
        test_data[2692] = 33'd2478811978;
        test_addr[2693] = 257;
        test_data[2693] = 33'd490540624;
        test_addr[2694] = 107;
        test_data[2694] = 33'd7661133238;
        test_addr[2695] = 835;
        test_data[2695] = 33'd135845962;
        test_addr[2696] = 625;
        test_data[2696] = 33'd8275388533;
        test_addr[2697] = 976;
        test_data[2697] = 33'd3395753456;
        test_addr[2698] = 810;
        test_data[2698] = 33'd3662887446;
        test_addr[2699] = 452;
        test_data[2699] = 33'd1875245374;
        test_addr[2700] = 177;
        test_data[2700] = 33'd2905827243;
        test_addr[2701] = 433;
        test_data[2701] = 33'd8519305820;
        test_addr[2702] = 334;
        test_data[2702] = 33'd6141804554;
        test_addr[2703] = 410;
        test_data[2703] = 33'd3670908267;
        test_addr[2704] = 489;
        test_data[2704] = 33'd4219814471;
        test_addr[2705] = 1016;
        test_data[2705] = 33'd5258863264;
        test_addr[2706] = 858;
        test_data[2706] = 33'd1864704728;
        test_addr[2707] = 745;
        test_data[2707] = 33'd5837527293;
        test_addr[2708] = 877;
        test_data[2708] = 33'd3606600498;
        test_addr[2709] = 962;
        test_data[2709] = 33'd1878395484;
        test_addr[2710] = 882;
        test_data[2710] = 33'd5953404875;
        test_addr[2711] = 308;
        test_data[2711] = 33'd5919315180;
        test_addr[2712] = 783;
        test_data[2712] = 33'd1379073191;
        test_addr[2713] = 558;
        test_data[2713] = 33'd6848915010;
        test_addr[2714] = 379;
        test_data[2714] = 33'd7144018043;
        test_addr[2715] = 337;
        test_data[2715] = 33'd3555484088;
        test_addr[2716] = 428;
        test_data[2716] = 33'd192890954;
        test_addr[2717] = 836;
        test_data[2717] = 33'd361379194;
        test_addr[2718] = 515;
        test_data[2718] = 33'd4537230457;
        test_addr[2719] = 597;
        test_data[2719] = 33'd2521741564;
        test_addr[2720] = 264;
        test_data[2720] = 33'd835312204;
        test_addr[2721] = 242;
        test_data[2721] = 33'd5485542569;
        test_addr[2722] = 29;
        test_data[2722] = 33'd1255285926;
        test_addr[2723] = 902;
        test_data[2723] = 33'd1242100171;
        test_addr[2724] = 52;
        test_data[2724] = 33'd5472781593;
        test_addr[2725] = 220;
        test_data[2725] = 33'd3833423383;
        test_addr[2726] = 717;
        test_data[2726] = 33'd2724895895;
        test_addr[2727] = 411;
        test_data[2727] = 33'd2424254182;
        test_addr[2728] = 176;
        test_data[2728] = 33'd799116268;
        test_addr[2729] = 115;
        test_data[2729] = 33'd4467948148;
        test_addr[2730] = 201;
        test_data[2730] = 33'd8393046847;
        test_addr[2731] = 657;
        test_data[2731] = 33'd8107453281;
        test_addr[2732] = 822;
        test_data[2732] = 33'd3946742381;
        test_addr[2733] = 852;
        test_data[2733] = 33'd3685315453;
        test_addr[2734] = 243;
        test_data[2734] = 33'd4020496137;
        test_addr[2735] = 1002;
        test_data[2735] = 33'd2359943401;
        test_addr[2736] = 850;
        test_data[2736] = 33'd2610616633;
        test_addr[2737] = 161;
        test_data[2737] = 33'd1596641998;
        test_addr[2738] = 331;
        test_data[2738] = 33'd2402963099;
        test_addr[2739] = 862;
        test_data[2739] = 33'd1299278838;
        test_addr[2740] = 85;
        test_data[2740] = 33'd6959272927;
        test_addr[2741] = 12;
        test_data[2741] = 33'd1981417174;
        test_addr[2742] = 769;
        test_data[2742] = 33'd5379517731;
        test_addr[2743] = 843;
        test_data[2743] = 33'd1336400027;
        test_addr[2744] = 839;
        test_data[2744] = 33'd5920045766;
        test_addr[2745] = 93;
        test_data[2745] = 33'd5878320782;
        test_addr[2746] = 449;
        test_data[2746] = 33'd2398926887;
        test_addr[2747] = 198;
        test_data[2747] = 33'd3924284121;
        test_addr[2748] = 335;
        test_data[2748] = 33'd3397286355;
        test_addr[2749] = 865;
        test_data[2749] = 33'd1670495772;
        test_addr[2750] = 299;
        test_data[2750] = 33'd3042141155;
        test_addr[2751] = 559;
        test_data[2751] = 33'd187816707;
        test_addr[2752] = 13;
        test_data[2752] = 33'd3216512318;
        test_addr[2753] = 626;
        test_data[2753] = 33'd132035543;
        test_addr[2754] = 384;
        test_data[2754] = 33'd547271751;
        test_addr[2755] = 779;
        test_data[2755] = 33'd4912899587;
        test_addr[2756] = 639;
        test_data[2756] = 33'd8112233422;
        test_addr[2757] = 644;
        test_data[2757] = 33'd2060679594;
        test_addr[2758] = 664;
        test_data[2758] = 33'd836176777;
        test_addr[2759] = 727;
        test_data[2759] = 33'd2548078876;
        test_addr[2760] = 466;
        test_data[2760] = 33'd7516324001;
        test_addr[2761] = 916;
        test_data[2761] = 33'd379022188;
        test_addr[2762] = 571;
        test_data[2762] = 33'd2554728556;
        test_addr[2763] = 336;
        test_data[2763] = 33'd5535498475;
        test_addr[2764] = 438;
        test_data[2764] = 33'd3272117358;
        test_addr[2765] = 653;
        test_data[2765] = 33'd3674868386;
        test_addr[2766] = 772;
        test_data[2766] = 33'd3207440178;
        test_addr[2767] = 631;
        test_data[2767] = 33'd1893022681;
        test_addr[2768] = 243;
        test_data[2768] = 33'd4020496137;
        test_addr[2769] = 505;
        test_data[2769] = 33'd3673032087;
        test_addr[2770] = 739;
        test_data[2770] = 33'd24113143;
        test_addr[2771] = 741;
        test_data[2771] = 33'd4313269272;
        test_addr[2772] = 765;
        test_data[2772] = 33'd843852261;
        test_addr[2773] = 617;
        test_data[2773] = 33'd306081816;
        test_addr[2774] = 728;
        test_data[2774] = 33'd2370403888;
        test_addr[2775] = 884;
        test_data[2775] = 33'd678817658;
        test_addr[2776] = 909;
        test_data[2776] = 33'd8408500060;
        test_addr[2777] = 974;
        test_data[2777] = 33'd7795562885;
        test_addr[2778] = 577;
        test_data[2778] = 33'd2874325634;
        test_addr[2779] = 11;
        test_data[2779] = 33'd5882696747;
        test_addr[2780] = 315;
        test_data[2780] = 33'd1859419918;
        test_addr[2781] = 414;
        test_data[2781] = 33'd4862343509;
        test_addr[2782] = 377;
        test_data[2782] = 33'd3153142852;
        test_addr[2783] = 150;
        test_data[2783] = 33'd4845491796;
        test_addr[2784] = 294;
        test_data[2784] = 33'd301140059;
        test_addr[2785] = 960;
        test_data[2785] = 33'd1617484150;
        test_addr[2786] = 625;
        test_data[2786] = 33'd3980421237;
        test_addr[2787] = 472;
        test_data[2787] = 33'd8383047452;
        test_addr[2788] = 288;
        test_data[2788] = 33'd262849900;
        test_addr[2789] = 1013;
        test_data[2789] = 33'd3443847325;
        test_addr[2790] = 727;
        test_data[2790] = 33'd2548078876;
        test_addr[2791] = 79;
        test_data[2791] = 33'd5861727944;
        test_addr[2792] = 640;
        test_data[2792] = 33'd2980138361;
        test_addr[2793] = 891;
        test_data[2793] = 33'd1858193830;
        test_addr[2794] = 245;
        test_data[2794] = 33'd1366539889;
        test_addr[2795] = 452;
        test_data[2795] = 33'd1875245374;
        test_addr[2796] = 161;
        test_data[2796] = 33'd1596641998;
        test_addr[2797] = 761;
        test_data[2797] = 33'd6210606249;
        test_addr[2798] = 375;
        test_data[2798] = 33'd796968996;
        test_addr[2799] = 893;
        test_data[2799] = 33'd3967042524;
        test_addr[2800] = 276;
        test_data[2800] = 33'd1049188557;
        test_addr[2801] = 556;
        test_data[2801] = 33'd1863958673;
        test_addr[2802] = 125;
        test_data[2802] = 33'd1259733705;
        test_addr[2803] = 70;
        test_data[2803] = 33'd5430648661;
        test_addr[2804] = 822;
        test_data[2804] = 33'd4813181398;
        test_addr[2805] = 116;
        test_data[2805] = 33'd6204490017;
        test_addr[2806] = 532;
        test_data[2806] = 33'd2499535484;
        test_addr[2807] = 579;
        test_data[2807] = 33'd2950567516;
        test_addr[2808] = 700;
        test_data[2808] = 33'd2118661662;
        test_addr[2809] = 169;
        test_data[2809] = 33'd6399581272;
        test_addr[2810] = 570;
        test_data[2810] = 33'd1605140899;
        test_addr[2811] = 955;
        test_data[2811] = 33'd1186627500;
        test_addr[2812] = 697;
        test_data[2812] = 33'd3895236155;
        test_addr[2813] = 1018;
        test_data[2813] = 33'd1157429103;
        test_addr[2814] = 50;
        test_data[2814] = 33'd1824887721;
        test_addr[2815] = 942;
        test_data[2815] = 33'd916379260;
        test_addr[2816] = 454;
        test_data[2816] = 33'd5673275776;
        test_addr[2817] = 696;
        test_data[2817] = 33'd3542107861;
        test_addr[2818] = 411;
        test_data[2818] = 33'd2424254182;
        test_addr[2819] = 34;
        test_data[2819] = 33'd5964364965;
        test_addr[2820] = 142;
        test_data[2820] = 33'd2263992737;
        test_addr[2821] = 185;
        test_data[2821] = 33'd804599567;
        test_addr[2822] = 1013;
        test_data[2822] = 33'd3443847325;
        test_addr[2823] = 865;
        test_data[2823] = 33'd1670495772;
        test_addr[2824] = 785;
        test_data[2824] = 33'd5048776861;
        test_addr[2825] = 356;
        test_data[2825] = 33'd5886822977;
        test_addr[2826] = 256;
        test_data[2826] = 33'd845636559;
        test_addr[2827] = 846;
        test_data[2827] = 33'd8463975280;
        test_addr[2828] = 659;
        test_data[2828] = 33'd3699990366;
        test_addr[2829] = 752;
        test_data[2829] = 33'd8245431519;
        test_addr[2830] = 78;
        test_data[2830] = 33'd6242519753;
        test_addr[2831] = 580;
        test_data[2831] = 33'd4090953264;
        test_addr[2832] = 240;
        test_data[2832] = 33'd4066667004;
        test_addr[2833] = 886;
        test_data[2833] = 33'd479387173;
        test_addr[2834] = 539;
        test_data[2834] = 33'd2220181209;
        test_addr[2835] = 620;
        test_data[2835] = 33'd990877164;
        test_addr[2836] = 292;
        test_data[2836] = 33'd1265860839;
        test_addr[2837] = 725;
        test_data[2837] = 33'd5543960032;
        test_addr[2838] = 335;
        test_data[2838] = 33'd3397286355;
        test_addr[2839] = 462;
        test_data[2839] = 33'd1029956024;
        test_addr[2840] = 705;
        test_data[2840] = 33'd4657010600;
        test_addr[2841] = 480;
        test_data[2841] = 33'd2118543923;
        test_addr[2842] = 697;
        test_data[2842] = 33'd3895236155;
        test_addr[2843] = 624;
        test_data[2843] = 33'd2766751231;
        test_addr[2844] = 773;
        test_data[2844] = 33'd531933772;
        test_addr[2845] = 851;
        test_data[2845] = 33'd852126570;
        test_addr[2846] = 895;
        test_data[2846] = 33'd3088967000;
        test_addr[2847] = 717;
        test_data[2847] = 33'd7457047552;
        test_addr[2848] = 666;
        test_data[2848] = 33'd3442547013;
        test_addr[2849] = 971;
        test_data[2849] = 33'd4477299893;
        test_addr[2850] = 959;
        test_data[2850] = 33'd88139643;
        test_addr[2851] = 394;
        test_data[2851] = 33'd2134209481;
        test_addr[2852] = 201;
        test_data[2852] = 33'd4098079551;
        test_addr[2853] = 717;
        test_data[2853] = 33'd3162080256;
        test_addr[2854] = 10;
        test_data[2854] = 33'd7750659633;
        test_addr[2855] = 603;
        test_data[2855] = 33'd2106932475;
        test_addr[2856] = 837;
        test_data[2856] = 33'd1693487156;
        test_addr[2857] = 192;
        test_data[2857] = 33'd740398394;
        test_addr[2858] = 570;
        test_data[2858] = 33'd1605140899;
        test_addr[2859] = 440;
        test_data[2859] = 33'd4898328579;
        test_addr[2860] = 976;
        test_data[2860] = 33'd7651203230;
        test_addr[2861] = 54;
        test_data[2861] = 33'd3762075597;
        test_addr[2862] = 834;
        test_data[2862] = 33'd2790802590;
        test_addr[2863] = 863;
        test_data[2863] = 33'd6879917381;
        test_addr[2864] = 532;
        test_data[2864] = 33'd8225515703;
        test_addr[2865] = 990;
        test_data[2865] = 33'd616895957;
        test_addr[2866] = 242;
        test_data[2866] = 33'd1190575273;
        test_addr[2867] = 699;
        test_data[2867] = 33'd3550875325;
        test_addr[2868] = 937;
        test_data[2868] = 33'd650004110;
        test_addr[2869] = 517;
        test_data[2869] = 33'd8473624721;
        test_addr[2870] = 223;
        test_data[2870] = 33'd3855190456;
        test_addr[2871] = 917;
        test_data[2871] = 33'd778607413;
        test_addr[2872] = 289;
        test_data[2872] = 33'd3920997515;
        test_addr[2873] = 0;
        test_data[2873] = 33'd3077293961;
        test_addr[2874] = 780;
        test_data[2874] = 33'd614300779;
        test_addr[2875] = 701;
        test_data[2875] = 33'd202904808;
        test_addr[2876] = 614;
        test_data[2876] = 33'd1386644667;
        test_addr[2877] = 1019;
        test_data[2877] = 33'd510091675;
        test_addr[2878] = 246;
        test_data[2878] = 33'd7864338706;
        test_addr[2879] = 565;
        test_data[2879] = 33'd4241384530;
        test_addr[2880] = 89;
        test_data[2880] = 33'd1425280291;
        test_addr[2881] = 864;
        test_data[2881] = 33'd4311950563;
        test_addr[2882] = 621;
        test_data[2882] = 33'd3667224622;
        test_addr[2883] = 163;
        test_data[2883] = 33'd3667441522;
        test_addr[2884] = 378;
        test_data[2884] = 33'd1591577112;
        test_addr[2885] = 173;
        test_data[2885] = 33'd285679836;
        test_addr[2886] = 409;
        test_data[2886] = 33'd1379904639;
        test_addr[2887] = 646;
        test_data[2887] = 33'd132734761;
        test_addr[2888] = 931;
        test_data[2888] = 33'd3388134606;
        test_addr[2889] = 87;
        test_data[2889] = 33'd3390580480;
        test_addr[2890] = 367;
        test_data[2890] = 33'd6764680167;
        test_addr[2891] = 731;
        test_data[2891] = 33'd6172711271;
        test_addr[2892] = 905;
        test_data[2892] = 33'd3962311491;
        test_addr[2893] = 241;
        test_data[2893] = 33'd1993840260;
        test_addr[2894] = 39;
        test_data[2894] = 33'd1662140024;
        test_addr[2895] = 978;
        test_data[2895] = 33'd1849704765;
        test_addr[2896] = 49;
        test_data[2896] = 33'd4201896278;
        test_addr[2897] = 91;
        test_data[2897] = 33'd961493540;
        test_addr[2898] = 583;
        test_data[2898] = 33'd5149294686;
        test_addr[2899] = 729;
        test_data[2899] = 33'd1893345796;
        test_addr[2900] = 842;
        test_data[2900] = 33'd7217382674;
        test_addr[2901] = 229;
        test_data[2901] = 33'd5823052937;
        test_addr[2902] = 399;
        test_data[2902] = 33'd2238490792;
        test_addr[2903] = 83;
        test_data[2903] = 33'd4027428377;
        test_addr[2904] = 17;
        test_data[2904] = 33'd567481263;
        test_addr[2905] = 571;
        test_data[2905] = 33'd2554728556;
        test_addr[2906] = 200;
        test_data[2906] = 33'd6345810720;
        test_addr[2907] = 457;
        test_data[2907] = 33'd4191839408;
        test_addr[2908] = 427;
        test_data[2908] = 33'd7166634916;
        test_addr[2909] = 346;
        test_data[2909] = 33'd355919171;
        test_addr[2910] = 678;
        test_data[2910] = 33'd3688685586;
        test_addr[2911] = 273;
        test_data[2911] = 33'd2277303350;
        test_addr[2912] = 100;
        test_data[2912] = 33'd5014102958;
        test_addr[2913] = 88;
        test_data[2913] = 33'd143353581;
        test_addr[2914] = 483;
        test_data[2914] = 33'd942928245;
        test_addr[2915] = 60;
        test_data[2915] = 33'd2293001596;
        test_addr[2916] = 847;
        test_data[2916] = 33'd4505703299;
        test_addr[2917] = 135;
        test_data[2917] = 33'd5909856631;
        test_addr[2918] = 97;
        test_data[2918] = 33'd62382029;
        test_addr[2919] = 888;
        test_data[2919] = 33'd685991554;
        test_addr[2920] = 636;
        test_data[2920] = 33'd5321758462;
        test_addr[2921] = 292;
        test_data[2921] = 33'd1265860839;
        test_addr[2922] = 945;
        test_data[2922] = 33'd1793343414;
        test_addr[2923] = 739;
        test_data[2923] = 33'd24113143;
        test_addr[2924] = 990;
        test_data[2924] = 33'd5376208957;
        test_addr[2925] = 906;
        test_data[2925] = 33'd4701813998;
        test_addr[2926] = 30;
        test_data[2926] = 33'd561337608;
        test_addr[2927] = 441;
        test_data[2927] = 33'd3607886437;
        test_addr[2928] = 767;
        test_data[2928] = 33'd1657730187;
        test_addr[2929] = 613;
        test_data[2929] = 33'd1975594517;
        test_addr[2930] = 609;
        test_data[2930] = 33'd779641857;
        test_addr[2931] = 197;
        test_data[2931] = 33'd4143794548;
        test_addr[2932] = 669;
        test_data[2932] = 33'd7662728341;
        test_addr[2933] = 386;
        test_data[2933] = 33'd4824001452;
        test_addr[2934] = 640;
        test_data[2934] = 33'd6495935681;
        test_addr[2935] = 465;
        test_data[2935] = 33'd4289052588;
        test_addr[2936] = 399;
        test_data[2936] = 33'd2238490792;
        test_addr[2937] = 535;
        test_data[2937] = 33'd553075824;
        test_addr[2938] = 129;
        test_data[2938] = 33'd3338914691;
        test_addr[2939] = 104;
        test_data[2939] = 33'd4499901015;
        test_addr[2940] = 341;
        test_data[2940] = 33'd720341552;
        test_addr[2941] = 107;
        test_data[2941] = 33'd3366165942;
        test_addr[2942] = 206;
        test_data[2942] = 33'd6380277275;
        test_addr[2943] = 970;
        test_data[2943] = 33'd8383159681;
        test_addr[2944] = 243;
        test_data[2944] = 33'd4020496137;
        test_addr[2945] = 114;
        test_data[2945] = 33'd5160014202;
        test_addr[2946] = 796;
        test_data[2946] = 33'd1296508384;
        test_addr[2947] = 151;
        test_data[2947] = 33'd6531236214;
        test_addr[2948] = 382;
        test_data[2948] = 33'd706838701;
        test_addr[2949] = 382;
        test_data[2949] = 33'd706838701;
        test_addr[2950] = 605;
        test_data[2950] = 33'd3854904784;
        test_addr[2951] = 1017;
        test_data[2951] = 33'd4360981718;
        test_addr[2952] = 34;
        test_data[2952] = 33'd1669397669;
        test_addr[2953] = 373;
        test_data[2953] = 33'd4092263069;
        test_addr[2954] = 641;
        test_data[2954] = 33'd2236541259;
        test_addr[2955] = 135;
        test_data[2955] = 33'd1614889335;
        test_addr[2956] = 510;
        test_data[2956] = 33'd195368792;
        test_addr[2957] = 185;
        test_data[2957] = 33'd804599567;
        test_addr[2958] = 203;
        test_data[2958] = 33'd6805699776;
        test_addr[2959] = 868;
        test_data[2959] = 33'd2145195459;
        test_addr[2960] = 740;
        test_data[2960] = 33'd5060931608;
        test_addr[2961] = 435;
        test_data[2961] = 33'd2086475014;
        test_addr[2962] = 324;
        test_data[2962] = 33'd1279699095;
        test_addr[2963] = 797;
        test_data[2963] = 33'd6581425702;
        test_addr[2964] = 489;
        test_data[2964] = 33'd4219814471;
        test_addr[2965] = 836;
        test_data[2965] = 33'd5294078423;
        test_addr[2966] = 913;
        test_data[2966] = 33'd803289427;
        test_addr[2967] = 714;
        test_data[2967] = 33'd5524770954;
        test_addr[2968] = 1014;
        test_data[2968] = 33'd8088898455;
        test_addr[2969] = 512;
        test_data[2969] = 33'd4210439056;
        test_addr[2970] = 945;
        test_data[2970] = 33'd1793343414;
        test_addr[2971] = 767;
        test_data[2971] = 33'd1657730187;
        test_addr[2972] = 901;
        test_data[2972] = 33'd2790845591;
        test_addr[2973] = 153;
        test_data[2973] = 33'd1670173968;
        test_addr[2974] = 901;
        test_data[2974] = 33'd2790845591;
        test_addr[2975] = 338;
        test_data[2975] = 33'd3638687009;
        test_addr[2976] = 537;
        test_data[2976] = 33'd1589033191;
        test_addr[2977] = 621;
        test_data[2977] = 33'd3667224622;
        test_addr[2978] = 588;
        test_data[2978] = 33'd4700321454;
        test_addr[2979] = 514;
        test_data[2979] = 33'd1348257185;
        test_addr[2980] = 525;
        test_data[2980] = 33'd4382258182;
        test_addr[2981] = 931;
        test_data[2981] = 33'd8131444315;
        test_addr[2982] = 78;
        test_data[2982] = 33'd1947552457;
        test_addr[2983] = 119;
        test_data[2983] = 33'd3348202238;
        test_addr[2984] = 451;
        test_data[2984] = 33'd2176493955;
        test_addr[2985] = 693;
        test_data[2985] = 33'd107943679;
        test_addr[2986] = 225;
        test_data[2986] = 33'd524980437;
        test_addr[2987] = 257;
        test_data[2987] = 33'd490540624;
        test_addr[2988] = 125;
        test_data[2988] = 33'd1259733705;
        test_addr[2989] = 858;
        test_data[2989] = 33'd8105707407;
        test_addr[2990] = 1015;
        test_data[2990] = 33'd4316194586;
        test_addr[2991] = 200;
        test_data[2991] = 33'd2050843424;
        test_addr[2992] = 578;
        test_data[2992] = 33'd5605780788;
        test_addr[2993] = 304;
        test_data[2993] = 33'd7902755669;
        test_addr[2994] = 483;
        test_data[2994] = 33'd6138281972;
        test_addr[2995] = 4;
        test_data[2995] = 33'd1143739882;
        test_addr[2996] = 567;
        test_data[2996] = 33'd4589564588;
        test_addr[2997] = 434;
        test_data[2997] = 33'd4825640152;
        test_addr[2998] = 188;
        test_data[2998] = 33'd1703939805;
        test_addr[2999] = 932;
        test_data[2999] = 33'd1842773940;

    end
endmodule
